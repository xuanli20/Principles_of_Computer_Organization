
/*
本文件是一个测试文件，用于测试cache模块
工作原理是模仿CPU的读写请求，对cache进行读写操作
将Cache返回的数据与预先数据进行比较，如果一致则测试通过
*/
`timescale 1ns/1ps
module cache_tb();

    //测试参数
    parameter READ_NUM = 2000;  // 测试次数 这里设置为2000次读，1000次写
    parameter WRITE_NUM = 1000;  
    //模块参数
    parameter INDEX_WIDTH       = 3;   // Cache索引位宽 2^3=8行
    parameter LINE_OFFSET_WIDTH = 2;   // 行偏移位宽，决定了一行的宽度 2^2=4字
    parameter SPACE_OFFSET      = 2;   // 一个地址空间占1个字节，因此一个字需要4个地址空间，由于假设为整字读取，处理地址的时候可以默认后两位为0
    parameter MEM_ADDR_WIDTH    = 10;   // 为了简化，这里假设内存地址宽度为10位（CPU请求地址仍然是32位，只不过我们这里简化处理，截断了高位） 
    parameter WAY_NUM           = 2;   // Cache N路组相联(N=1的时候是直接映射)

    // 变化的信号 CPU发出
    reg clk=1;
    reg rstn=1;
    reg stat=0;
    // 等rstn信号稳定后 clk信号才开始翻转
    initial begin
        #1 rstn = 0;
        #1 rstn = 1;
        stat = 1;
    end
    always  #1 clk = ~clk;

    wire [31:0] addr;
    wire r_req;
    wire w_req;
    wire [31:0] w_data;

    // 导线
    wire [31:0] r_data;
    wire miss;
    wire mem_r;
    wire mem_w;
    wire [31:0] mem_addr;
    wire [127:0] mem_w_data;
    wire [127:0] mem_r_data;
    wire mem_ready;

    // 用于测试的信号
    reg [MEM_ADDR_WIDTH-1:0] test_addr[0:READ_NUM+WRITE_NUM-1];  // 用于存储测试地址
    reg [32:0] test_data[0:READ_NUM+WRITE_NUM-1];  // 用于存储测试数据 最高位用于标记是否写入 0：读 1：写
    reg [31:0] test_cnt=0;  // 用于计数，每次读写操作后加1
    reg diff=0;  // 用于标记是否有不一致的数据

    // 用于对比的提交，当前cache应该给出的数据
    wire op;
    wire[31:0] data;
    assign op = test_data[test_cnt-1][32];
    assign data = test_data[test_cnt-1][31:0];
    
    // 状态机
    assign addr = test_addr[test_cnt]<<SPACE_OFFSET;
    assign r_req = test_data[test_cnt][32] == 0 ? 1 : 0;
    assign w_req = test_data[test_cnt][32] == 1 ? 1 : 0;
    assign w_data = test_data[test_cnt][31:0];
    always @(posedge clk) begin
        if (!miss && (test_cnt < READ_NUM+WRITE_NUM) && stat) begin
            if (test_data[test_cnt-1][32] == 0) begin  // 读
                if (r_data != test_data[test_cnt-1][31:0]) begin
                    $display("Read error at %d, expect %h, get %h", test_cnt, test_data[test_cnt-1][31:0], r_data);
                    diff = 1;
                end
            end
            test_cnt <= test_cnt + 1;
        end
    end

    // 例化cache
    cache_random #(
        .INDEX_WIDTH(INDEX_WIDTH),
        .LINE_OFFSET_WIDTH(LINE_OFFSET_WIDTH),
        .SPACE_OFFSET(SPACE_OFFSET),
        .WAY_NUM(WAY_NUM),
        .N(1)
    ) cache(
        .clk(clk),
        .rstn(rstn),
        .addr(addr),
        .r_req(r_req),
        .w_req(w_req),
        .w_data(w_data),
        .r_data(r_data),
        .miss(miss),
        .mem_r(mem_r),
        .mem_w(mem_w),
        .mem_addr(mem_addr),
        .mem_w_data(mem_w_data),
        .mem_r_data(mem_r_data),
        .mem_ready(mem_ready)
    );

    // 内存
    mem #(
        .INDEX_WIDTH(INDEX_WIDTH),
        .LINE_OFFSET_WIDTH(LINE_OFFSET_WIDTH),
        .SPACE_OFFSET(SPACE_OFFSET),
        .MEM_ADDR_WIDTH(MEM_ADDR_WIDTH-LINE_OFFSET_WIDTH),
        .WAY_NUM(WAY_NUM)
    ) mem_inst(
        .clk(clk),
        .rstn(rstn),
        .mem_r(mem_r),
        .mem_w(mem_w),
        .mem_addr(mem_addr),
        .mem_w_data(mem_w_data),
        .mem_r_data(mem_r_data),
        .mem_ready(mem_ready)
    );

    // 初始化测试数据
    initial begin
        test_addr[0] = 0;
        test_data[0] = 33'd812361294;
        test_addr[1] = 1;
        test_data[1] = 33'd1897396466;
        test_addr[2] = 2;
        test_data[2] = 33'd6160420735;
        test_addr[3] = 3;
        test_data[3] = 33'd5306660553;
        test_addr[4] = 4;
        test_data[4] = 33'd4388524592;
        test_addr[5] = 527;
        test_data[5] = 33'd3681101907;
        test_addr[6] = 528;
        test_data[6] = 33'd1983832739;
        test_addr[7] = 529;
        test_data[7] = 33'd3177420342;
        test_addr[8] = 530;
        test_data[8] = 33'd7328527154;
        test_addr[9] = 531;
        test_data[9] = 33'd4269338406;
        test_addr[10] = 532;
        test_data[10] = 33'd1758387349;
        test_addr[11] = 533;
        test_data[11] = 33'd3892039782;
        test_addr[12] = 534;
        test_data[12] = 33'd3083492837;
        test_addr[13] = 535;
        test_data[13] = 33'd4630439284;
        test_addr[14] = 536;
        test_data[14] = 33'd3377477922;
        test_addr[15] = 537;
        test_data[15] = 33'd1309125160;
        test_addr[16] = 538;
        test_data[16] = 33'd1250172866;
        test_addr[17] = 539;
        test_data[17] = 33'd6633252007;
        test_addr[18] = 540;
        test_data[18] = 33'd5660260884;
        test_addr[19] = 541;
        test_data[19] = 33'd3682747475;
        test_addr[20] = 5;
        test_data[20] = 33'd5723413021;
        test_addr[21] = 6;
        test_data[21] = 33'd1309544095;
        test_addr[22] = 7;
        test_data[22] = 33'd3491080214;
        test_addr[23] = 460;
        test_data[23] = 33'd2977339794;
        test_addr[24] = 8;
        test_data[24] = 33'd1793239769;
        test_addr[25] = 9;
        test_data[25] = 33'd1174159001;
        test_addr[26] = 699;
        test_data[26] = 33'd7975476024;
        test_addr[27] = 700;
        test_data[27] = 33'd5648057908;
        test_addr[28] = 701;
        test_data[28] = 33'd3933897631;
        test_addr[29] = 702;
        test_data[29] = 33'd6196517671;
        test_addr[30] = 10;
        test_data[30] = 33'd1664182063;
        test_addr[31] = 11;
        test_data[31] = 33'd773081521;
        test_addr[32] = 12;
        test_data[32] = 33'd3296343955;
        test_addr[33] = 13;
        test_data[33] = 33'd1476987912;
        test_addr[34] = 14;
        test_data[34] = 33'd1747019271;
        test_addr[35] = 15;
        test_data[35] = 33'd5684875099;
        test_addr[36] = 16;
        test_data[36] = 33'd7290688680;
        test_addr[37] = 17;
        test_data[37] = 33'd1707974702;
        test_addr[38] = 18;
        test_data[38] = 33'd5866918601;
        test_addr[39] = 19;
        test_data[39] = 33'd1943724055;
        test_addr[40] = 20;
        test_data[40] = 33'd1223440380;
        test_addr[41] = 21;
        test_data[41] = 33'd3366782182;
        test_addr[42] = 22;
        test_data[42] = 33'd883716006;
        test_addr[43] = 23;
        test_data[43] = 33'd2361297799;
        test_addr[44] = 24;
        test_data[44] = 33'd2711593210;
        test_addr[45] = 25;
        test_data[45] = 33'd4002336428;
        test_addr[46] = 26;
        test_data[46] = 33'd4291600053;
        test_addr[47] = 27;
        test_data[47] = 33'd4539737994;
        test_addr[48] = 28;
        test_data[48] = 33'd1899814066;
        test_addr[49] = 29;
        test_data[49] = 33'd3331445440;
        test_addr[50] = 30;
        test_data[50] = 33'd1741498846;
        test_addr[51] = 31;
        test_data[51] = 33'd4308069556;
        test_addr[52] = 32;
        test_data[52] = 33'd1170076186;
        test_addr[53] = 33;
        test_data[53] = 33'd2359621732;
        test_addr[54] = 34;
        test_data[54] = 33'd1887051034;
        test_addr[55] = 35;
        test_data[55] = 33'd4467650907;
        test_addr[56] = 36;
        test_data[56] = 33'd2709550290;
        test_addr[57] = 37;
        test_data[57] = 33'd406326701;
        test_addr[58] = 38;
        test_data[58] = 33'd3133901872;
        test_addr[59] = 39;
        test_data[59] = 33'd1715945728;
        test_addr[60] = 40;
        test_data[60] = 33'd3642725099;
        test_addr[61] = 41;
        test_data[61] = 33'd2411058451;
        test_addr[62] = 42;
        test_data[62] = 33'd7154381702;
        test_addr[63] = 43;
        test_data[63] = 33'd389770497;
        test_addr[64] = 44;
        test_data[64] = 33'd2890247156;
        test_addr[65] = 45;
        test_data[65] = 33'd1444532856;
        test_addr[66] = 46;
        test_data[66] = 33'd2921447489;
        test_addr[67] = 47;
        test_data[67] = 33'd6979472559;
        test_addr[68] = 48;
        test_data[68] = 33'd64235302;
        test_addr[69] = 49;
        test_data[69] = 33'd1390656163;
        test_addr[70] = 50;
        test_data[70] = 33'd2480296893;
        test_addr[71] = 573;
        test_data[71] = 33'd4029761842;
        test_addr[72] = 51;
        test_data[72] = 33'd893530107;
        test_addr[73] = 52;
        test_data[73] = 33'd369651485;
        test_addr[74] = 53;
        test_data[74] = 33'd2187729913;
        test_addr[75] = 54;
        test_data[75] = 33'd1681690332;
        test_addr[76] = 55;
        test_data[76] = 33'd1478733057;
        test_addr[77] = 56;
        test_data[77] = 33'd13033719;
        test_addr[78] = 57;
        test_data[78] = 33'd7780685032;
        test_addr[79] = 58;
        test_data[79] = 33'd528146972;
        test_addr[80] = 59;
        test_data[80] = 33'd7787481827;
        test_addr[81] = 60;
        test_data[81] = 33'd2587167315;
        test_addr[82] = 61;
        test_data[82] = 33'd3444518270;
        test_addr[83] = 62;
        test_data[83] = 33'd2627318154;
        test_addr[84] = 63;
        test_data[84] = 33'd12778738;
        test_addr[85] = 64;
        test_data[85] = 33'd4280548596;
        test_addr[86] = 978;
        test_data[86] = 33'd5817144597;
        test_addr[87] = 979;
        test_data[87] = 33'd3351282188;
        test_addr[88] = 980;
        test_data[88] = 33'd127768736;
        test_addr[89] = 981;
        test_data[89] = 33'd8173223286;
        test_addr[90] = 982;
        test_data[90] = 33'd5677731019;
        test_addr[91] = 983;
        test_data[91] = 33'd1650122225;
        test_addr[92] = 65;
        test_data[92] = 33'd3000665519;
        test_addr[93] = 208;
        test_data[93] = 33'd6522065189;
        test_addr[94] = 209;
        test_data[94] = 33'd7961997028;
        test_addr[95] = 210;
        test_data[95] = 33'd2312377961;
        test_addr[96] = 211;
        test_data[96] = 33'd2875926310;
        test_addr[97] = 212;
        test_data[97] = 33'd2392747211;
        test_addr[98] = 213;
        test_data[98] = 33'd7254391394;
        test_addr[99] = 214;
        test_data[99] = 33'd7365694971;
        test_addr[100] = 215;
        test_data[100] = 33'd7249970957;
        test_addr[101] = 216;
        test_data[101] = 33'd2609755010;
        test_addr[102] = 217;
        test_data[102] = 33'd1119239002;
        test_addr[103] = 218;
        test_data[103] = 33'd2296008684;
        test_addr[104] = 219;
        test_data[104] = 33'd3225055293;
        test_addr[105] = 220;
        test_data[105] = 33'd5966289262;
        test_addr[106] = 221;
        test_data[106] = 33'd1801818893;
        test_addr[107] = 222;
        test_data[107] = 33'd727510908;
        test_addr[108] = 223;
        test_data[108] = 33'd2764688405;
        test_addr[109] = 224;
        test_data[109] = 33'd6621989380;
        test_addr[110] = 225;
        test_data[110] = 33'd3019194714;
        test_addr[111] = 226;
        test_data[111] = 33'd8576816678;
        test_addr[112] = 227;
        test_data[112] = 33'd1667423717;
        test_addr[113] = 228;
        test_data[113] = 33'd1082603118;
        test_addr[114] = 229;
        test_data[114] = 33'd1506219133;
        test_addr[115] = 230;
        test_data[115] = 33'd3332009274;
        test_addr[116] = 66;
        test_data[116] = 33'd2358437066;
        test_addr[117] = 67;
        test_data[117] = 33'd1974385293;
        test_addr[118] = 68;
        test_data[118] = 33'd1457236560;
        test_addr[119] = 69;
        test_data[119] = 33'd912614945;
        test_addr[120] = 586;
        test_data[120] = 33'd3407577517;
        test_addr[121] = 587;
        test_data[121] = 33'd976124543;
        test_addr[122] = 588;
        test_data[122] = 33'd1568993292;
        test_addr[123] = 589;
        test_data[123] = 33'd1522418319;
        test_addr[124] = 590;
        test_data[124] = 33'd3186803448;
        test_addr[125] = 591;
        test_data[125] = 33'd5015581341;
        test_addr[126] = 70;
        test_data[126] = 33'd4479801324;
        test_addr[127] = 869;
        test_data[127] = 33'd6345471904;
        test_addr[128] = 870;
        test_data[128] = 33'd2235229089;
        test_addr[129] = 871;
        test_data[129] = 33'd3307625235;
        test_addr[130] = 872;
        test_data[130] = 33'd7793902835;
        test_addr[131] = 873;
        test_data[131] = 33'd7078549127;
        test_addr[132] = 874;
        test_data[132] = 33'd3793369460;
        test_addr[133] = 875;
        test_data[133] = 33'd4043269648;
        test_addr[134] = 876;
        test_data[134] = 33'd1362121102;
        test_addr[135] = 877;
        test_data[135] = 33'd2198385985;
        test_addr[136] = 878;
        test_data[136] = 33'd886953612;
        test_addr[137] = 879;
        test_data[137] = 33'd3146529035;
        test_addr[138] = 71;
        test_data[138] = 33'd7210879693;
        test_addr[139] = 72;
        test_data[139] = 33'd5751059807;
        test_addr[140] = 73;
        test_data[140] = 33'd3301388465;
        test_addr[141] = 74;
        test_data[141] = 33'd2014563986;
        test_addr[142] = 75;
        test_data[142] = 33'd7101044940;
        test_addr[143] = 76;
        test_data[143] = 33'd6737920874;
        test_addr[144] = 77;
        test_data[144] = 33'd7257034855;
        test_addr[145] = 78;
        test_data[145] = 33'd6520410432;
        test_addr[146] = 826;
        test_data[146] = 33'd251042263;
        test_addr[147] = 79;
        test_data[147] = 33'd1775955632;
        test_addr[148] = 80;
        test_data[148] = 33'd8022711996;
        test_addr[149] = 81;
        test_data[149] = 33'd3550050089;
        test_addr[150] = 82;
        test_data[150] = 33'd1564001926;
        test_addr[151] = 83;
        test_data[151] = 33'd1729932993;
        test_addr[152] = 84;
        test_data[152] = 33'd8256787361;
        test_addr[153] = 85;
        test_data[153] = 33'd2686387223;
        test_addr[154] = 86;
        test_data[154] = 33'd6046932994;
        test_addr[155] = 87;
        test_data[155] = 33'd5442979426;
        test_addr[156] = 88;
        test_data[156] = 33'd2879312064;
        test_addr[157] = 89;
        test_data[157] = 33'd8226503311;
        test_addr[158] = 90;
        test_data[158] = 33'd3551737466;
        test_addr[159] = 91;
        test_data[159] = 33'd1285586415;
        test_addr[160] = 92;
        test_data[160] = 33'd7041548576;
        test_addr[161] = 93;
        test_data[161] = 33'd8055773630;
        test_addr[162] = 94;
        test_data[162] = 33'd2987649344;
        test_addr[163] = 95;
        test_data[163] = 33'd2737991781;
        test_addr[164] = 96;
        test_data[164] = 33'd3739168123;
        test_addr[165] = 97;
        test_data[165] = 33'd1649687892;
        test_addr[166] = 98;
        test_data[166] = 33'd5437313110;
        test_addr[167] = 99;
        test_data[167] = 33'd3659483916;
        test_addr[168] = 100;
        test_data[168] = 33'd1882137235;
        test_addr[169] = 101;
        test_data[169] = 33'd7284935600;
        test_addr[170] = 836;
        test_data[170] = 33'd2037704408;
        test_addr[171] = 837;
        test_data[171] = 33'd1657911559;
        test_addr[172] = 838;
        test_data[172] = 33'd924586107;
        test_addr[173] = 839;
        test_data[173] = 33'd1862425237;
        test_addr[174] = 840;
        test_data[174] = 33'd8585264598;
        test_addr[175] = 841;
        test_data[175] = 33'd209372675;
        test_addr[176] = 842;
        test_data[176] = 33'd2607202746;
        test_addr[177] = 843;
        test_data[177] = 33'd4105319985;
        test_addr[178] = 844;
        test_data[178] = 33'd4108930760;
        test_addr[179] = 845;
        test_data[179] = 33'd3010963361;
        test_addr[180] = 846;
        test_data[180] = 33'd3871268654;
        test_addr[181] = 847;
        test_data[181] = 33'd2811533726;
        test_addr[182] = 848;
        test_data[182] = 33'd6284115384;
        test_addr[183] = 849;
        test_data[183] = 33'd4029825875;
        test_addr[184] = 850;
        test_data[184] = 33'd8154437474;
        test_addr[185] = 851;
        test_data[185] = 33'd3497740514;
        test_addr[186] = 852;
        test_data[186] = 33'd2241971371;
        test_addr[187] = 853;
        test_data[187] = 33'd2928255153;
        test_addr[188] = 854;
        test_data[188] = 33'd8547341066;
        test_addr[189] = 855;
        test_data[189] = 33'd2688237503;
        test_addr[190] = 856;
        test_data[190] = 33'd3274644583;
        test_addr[191] = 857;
        test_data[191] = 33'd2231454879;
        test_addr[192] = 858;
        test_data[192] = 33'd4000613725;
        test_addr[193] = 859;
        test_data[193] = 33'd544317971;
        test_addr[194] = 860;
        test_data[194] = 33'd3246602886;
        test_addr[195] = 861;
        test_data[195] = 33'd1495467381;
        test_addr[196] = 862;
        test_data[196] = 33'd3532219985;
        test_addr[197] = 863;
        test_data[197] = 33'd2533925369;
        test_addr[198] = 864;
        test_data[198] = 33'd5074511919;
        test_addr[199] = 865;
        test_data[199] = 33'd3491167284;
        test_addr[200] = 866;
        test_data[200] = 33'd4579011847;
        test_addr[201] = 867;
        test_data[201] = 33'd4306595764;
        test_addr[202] = 868;
        test_data[202] = 33'd3743578642;
        test_addr[203] = 869;
        test_data[203] = 33'd2050504608;
        test_addr[204] = 870;
        test_data[204] = 33'd2235229089;
        test_addr[205] = 102;
        test_data[205] = 33'd8068095491;
        test_addr[206] = 103;
        test_data[206] = 33'd1019640399;
        test_addr[207] = 104;
        test_data[207] = 33'd5616851972;
        test_addr[208] = 105;
        test_data[208] = 33'd627517218;
        test_addr[209] = 106;
        test_data[209] = 33'd5261072462;
        test_addr[210] = 107;
        test_data[210] = 33'd3217439098;
        test_addr[211] = 108;
        test_data[211] = 33'd8031918274;
        test_addr[212] = 109;
        test_data[212] = 33'd264822472;
        test_addr[213] = 110;
        test_data[213] = 33'd4027024129;
        test_addr[214] = 111;
        test_data[214] = 33'd645329535;
        test_addr[215] = 112;
        test_data[215] = 33'd6110608750;
        test_addr[216] = 113;
        test_data[216] = 33'd4144529833;
        test_addr[217] = 114;
        test_data[217] = 33'd2554819996;
        test_addr[218] = 115;
        test_data[218] = 33'd3969435406;
        test_addr[219] = 116;
        test_data[219] = 33'd1512917393;
        test_addr[220] = 117;
        test_data[220] = 33'd3459749905;
        test_addr[221] = 118;
        test_data[221] = 33'd2078089603;
        test_addr[222] = 747;
        test_data[222] = 33'd7510016708;
        test_addr[223] = 748;
        test_data[223] = 33'd8130941222;
        test_addr[224] = 749;
        test_data[224] = 33'd3249465326;
        test_addr[225] = 750;
        test_data[225] = 33'd3873234694;
        test_addr[226] = 751;
        test_data[226] = 33'd2207759834;
        test_addr[227] = 752;
        test_data[227] = 33'd5686836075;
        test_addr[228] = 753;
        test_data[228] = 33'd5076807933;
        test_addr[229] = 754;
        test_data[229] = 33'd7529714689;
        test_addr[230] = 755;
        test_data[230] = 33'd2779572929;
        test_addr[231] = 119;
        test_data[231] = 33'd5618322396;
        test_addr[232] = 120;
        test_data[232] = 33'd557041591;
        test_addr[233] = 121;
        test_data[233] = 33'd4852146673;
        test_addr[234] = 122;
        test_data[234] = 33'd886188703;
        test_addr[235] = 123;
        test_data[235] = 33'd978523342;
        test_addr[236] = 124;
        test_data[236] = 33'd2261534157;
        test_addr[237] = 125;
        test_data[237] = 33'd4331761732;
        test_addr[238] = 126;
        test_data[238] = 33'd717632510;
        test_addr[239] = 127;
        test_data[239] = 33'd6131785932;
        test_addr[240] = 128;
        test_data[240] = 33'd8380543487;
        test_addr[241] = 129;
        test_data[241] = 33'd438601362;
        test_addr[242] = 130;
        test_data[242] = 33'd2760717433;
        test_addr[243] = 131;
        test_data[243] = 33'd3219734873;
        test_addr[244] = 132;
        test_data[244] = 33'd1457531679;
        test_addr[245] = 133;
        test_data[245] = 33'd5460120569;
        test_addr[246] = 134;
        test_data[246] = 33'd7791061935;
        test_addr[247] = 135;
        test_data[247] = 33'd3470509274;
        test_addr[248] = 136;
        test_data[248] = 33'd5661493515;
        test_addr[249] = 137;
        test_data[249] = 33'd4277997269;
        test_addr[250] = 138;
        test_data[250] = 33'd51940499;
        test_addr[251] = 139;
        test_data[251] = 33'd4250352825;
        test_addr[252] = 512;
        test_data[252] = 33'd8187029204;
        test_addr[253] = 513;
        test_data[253] = 33'd45075662;
        test_addr[254] = 514;
        test_data[254] = 33'd8103272599;
        test_addr[255] = 515;
        test_data[255] = 33'd934899158;
        test_addr[256] = 516;
        test_data[256] = 33'd6203025336;
        test_addr[257] = 517;
        test_data[257] = 33'd1106079426;
        test_addr[258] = 518;
        test_data[258] = 33'd209533787;
        test_addr[259] = 519;
        test_data[259] = 33'd2029500360;
        test_addr[260] = 520;
        test_data[260] = 33'd6149215146;
        test_addr[261] = 521;
        test_data[261] = 33'd1928735641;
        test_addr[262] = 522;
        test_data[262] = 33'd6254841440;
        test_addr[263] = 523;
        test_data[263] = 33'd3215894844;
        test_addr[264] = 524;
        test_data[264] = 33'd3814837793;
        test_addr[265] = 525;
        test_data[265] = 33'd7263803437;
        test_addr[266] = 140;
        test_data[266] = 33'd4859584815;
        test_addr[267] = 141;
        test_data[267] = 33'd485567310;
        test_addr[268] = 142;
        test_data[268] = 33'd1458947625;
        test_addr[269] = 143;
        test_data[269] = 33'd730436975;
        test_addr[270] = 272;
        test_data[270] = 33'd3539921614;
        test_addr[271] = 273;
        test_data[271] = 33'd7986966442;
        test_addr[272] = 144;
        test_data[272] = 33'd7950431324;
        test_addr[273] = 145;
        test_data[273] = 33'd5311470609;
        test_addr[274] = 146;
        test_data[274] = 33'd1483917544;
        test_addr[275] = 147;
        test_data[275] = 33'd3933851125;
        test_addr[276] = 148;
        test_data[276] = 33'd1074274996;
        test_addr[277] = 149;
        test_data[277] = 33'd304283732;
        test_addr[278] = 150;
        test_data[278] = 33'd1383869392;
        test_addr[279] = 151;
        test_data[279] = 33'd2820628440;
        test_addr[280] = 152;
        test_data[280] = 33'd5621878822;
        test_addr[281] = 153;
        test_data[281] = 33'd327985978;
        test_addr[282] = 154;
        test_data[282] = 33'd412214464;
        test_addr[283] = 155;
        test_data[283] = 33'd3182442945;
        test_addr[284] = 5;
        test_data[284] = 33'd5133654741;
        test_addr[285] = 6;
        test_data[285] = 33'd7569268206;
        test_addr[286] = 156;
        test_data[286] = 33'd4176867573;
        test_addr[287] = 157;
        test_data[287] = 33'd1333860272;
        test_addr[288] = 158;
        test_data[288] = 33'd4087206092;
        test_addr[289] = 159;
        test_data[289] = 33'd7223563233;
        test_addr[290] = 160;
        test_data[290] = 33'd4955884555;
        test_addr[291] = 161;
        test_data[291] = 33'd8119335094;
        test_addr[292] = 162;
        test_data[292] = 33'd1461900145;
        test_addr[293] = 163;
        test_data[293] = 33'd6629793676;
        test_addr[294] = 164;
        test_data[294] = 33'd617221806;
        test_addr[295] = 165;
        test_data[295] = 33'd117310100;
        test_addr[296] = 166;
        test_data[296] = 33'd2648221725;
        test_addr[297] = 167;
        test_data[297] = 33'd7936482672;
        test_addr[298] = 168;
        test_data[298] = 33'd254554983;
        test_addr[299] = 169;
        test_data[299] = 33'd5859729520;
        test_addr[300] = 170;
        test_data[300] = 33'd574793399;
        test_addr[301] = 171;
        test_data[301] = 33'd753209148;
        test_addr[302] = 172;
        test_data[302] = 33'd460255681;
        test_addr[303] = 173;
        test_data[303] = 33'd5333902921;
        test_addr[304] = 174;
        test_data[304] = 33'd1373713971;
        test_addr[305] = 175;
        test_data[305] = 33'd5316358621;
        test_addr[306] = 176;
        test_data[306] = 33'd2743796502;
        test_addr[307] = 177;
        test_data[307] = 33'd1825087556;
        test_addr[308] = 178;
        test_data[308] = 33'd3775849174;
        test_addr[309] = 179;
        test_data[309] = 33'd1928357839;
        test_addr[310] = 236;
        test_data[310] = 33'd7307377236;
        test_addr[311] = 237;
        test_data[311] = 33'd168920287;
        test_addr[312] = 238;
        test_data[312] = 33'd4682825458;
        test_addr[313] = 239;
        test_data[313] = 33'd3601678559;
        test_addr[314] = 240;
        test_data[314] = 33'd4567368956;
        test_addr[315] = 241;
        test_data[315] = 33'd1202615656;
        test_addr[316] = 242;
        test_data[316] = 33'd1167664452;
        test_addr[317] = 243;
        test_data[317] = 33'd6299246270;
        test_addr[318] = 244;
        test_data[318] = 33'd1146573824;
        test_addr[319] = 245;
        test_data[319] = 33'd4434282718;
        test_addr[320] = 246;
        test_data[320] = 33'd4643287289;
        test_addr[321] = 247;
        test_data[321] = 33'd5533670862;
        test_addr[322] = 248;
        test_data[322] = 33'd7836453525;
        test_addr[323] = 249;
        test_data[323] = 33'd230942795;
        test_addr[324] = 250;
        test_data[324] = 33'd157822933;
        test_addr[325] = 251;
        test_data[325] = 33'd2172745435;
        test_addr[326] = 252;
        test_data[326] = 33'd3216848485;
        test_addr[327] = 253;
        test_data[327] = 33'd522192966;
        test_addr[328] = 254;
        test_data[328] = 33'd4309304770;
        test_addr[329] = 255;
        test_data[329] = 33'd714439378;
        test_addr[330] = 256;
        test_data[330] = 33'd2800244347;
        test_addr[331] = 257;
        test_data[331] = 33'd248550902;
        test_addr[332] = 258;
        test_data[332] = 33'd8171881359;
        test_addr[333] = 259;
        test_data[333] = 33'd2756113887;
        test_addr[334] = 260;
        test_data[334] = 33'd1766135903;
        test_addr[335] = 261;
        test_data[335] = 33'd4204582623;
        test_addr[336] = 180;
        test_data[336] = 33'd3962182398;
        test_addr[337] = 181;
        test_data[337] = 33'd5790772110;
        test_addr[338] = 182;
        test_data[338] = 33'd557477877;
        test_addr[339] = 183;
        test_data[339] = 33'd1320690480;
        test_addr[340] = 184;
        test_data[340] = 33'd7502115262;
        test_addr[341] = 185;
        test_data[341] = 33'd76388760;
        test_addr[342] = 186;
        test_data[342] = 33'd3665623001;
        test_addr[343] = 187;
        test_data[343] = 33'd800185981;
        test_addr[344] = 188;
        test_data[344] = 33'd7812163549;
        test_addr[345] = 189;
        test_data[345] = 33'd3256549792;
        test_addr[346] = 190;
        test_data[346] = 33'd6668816859;
        test_addr[347] = 191;
        test_data[347] = 33'd7029035031;
        test_addr[348] = 192;
        test_data[348] = 33'd5711076665;
        test_addr[349] = 193;
        test_data[349] = 33'd6958456400;
        test_addr[350] = 194;
        test_data[350] = 33'd117118296;
        test_addr[351] = 451;
        test_data[351] = 33'd8238727371;
        test_addr[352] = 452;
        test_data[352] = 33'd4299775126;
        test_addr[353] = 453;
        test_data[353] = 33'd1872832286;
        test_addr[354] = 454;
        test_data[354] = 33'd6414796394;
        test_addr[355] = 455;
        test_data[355] = 33'd2792297812;
        test_addr[356] = 456;
        test_data[356] = 33'd7006142339;
        test_addr[357] = 195;
        test_data[357] = 33'd4579747108;
        test_addr[358] = 196;
        test_data[358] = 33'd1622317500;
        test_addr[359] = 197;
        test_data[359] = 33'd2750204444;
        test_addr[360] = 198;
        test_data[360] = 33'd4651466781;
        test_addr[361] = 648;
        test_data[361] = 33'd776883759;
        test_addr[362] = 649;
        test_data[362] = 33'd3154846827;
        test_addr[363] = 650;
        test_data[363] = 33'd1968337716;
        test_addr[364] = 651;
        test_data[364] = 33'd7061204518;
        test_addr[365] = 652;
        test_data[365] = 33'd1737322648;
        test_addr[366] = 653;
        test_data[366] = 33'd7653683482;
        test_addr[367] = 654;
        test_data[367] = 33'd6249999459;
        test_addr[368] = 655;
        test_data[368] = 33'd3509997369;
        test_addr[369] = 656;
        test_data[369] = 33'd218457727;
        test_addr[370] = 657;
        test_data[370] = 33'd8368605320;
        test_addr[371] = 658;
        test_data[371] = 33'd420911824;
        test_addr[372] = 659;
        test_data[372] = 33'd3715143865;
        test_addr[373] = 660;
        test_data[373] = 33'd270341019;
        test_addr[374] = 661;
        test_data[374] = 33'd3720845072;
        test_addr[375] = 662;
        test_data[375] = 33'd2741441705;
        test_addr[376] = 663;
        test_data[376] = 33'd2417445093;
        test_addr[377] = 664;
        test_data[377] = 33'd961409848;
        test_addr[378] = 665;
        test_data[378] = 33'd7732823185;
        test_addr[379] = 666;
        test_data[379] = 33'd3656350260;
        test_addr[380] = 667;
        test_data[380] = 33'd6453846923;
        test_addr[381] = 668;
        test_data[381] = 33'd6641148744;
        test_addr[382] = 669;
        test_data[382] = 33'd420503772;
        test_addr[383] = 670;
        test_data[383] = 33'd2483701347;
        test_addr[384] = 671;
        test_data[384] = 33'd660543359;
        test_addr[385] = 672;
        test_data[385] = 33'd7952311023;
        test_addr[386] = 673;
        test_data[386] = 33'd3460743945;
        test_addr[387] = 674;
        test_data[387] = 33'd1495437377;
        test_addr[388] = 675;
        test_data[388] = 33'd3828766155;
        test_addr[389] = 676;
        test_data[389] = 33'd1442188537;
        test_addr[390] = 677;
        test_data[390] = 33'd4176733826;
        test_addr[391] = 678;
        test_data[391] = 33'd7270806388;
        test_addr[392] = 679;
        test_data[392] = 33'd1411385993;
        test_addr[393] = 680;
        test_data[393] = 33'd8156931980;
        test_addr[394] = 681;
        test_data[394] = 33'd7665304350;
        test_addr[395] = 682;
        test_data[395] = 33'd4475182272;
        test_addr[396] = 683;
        test_data[396] = 33'd452619150;
        test_addr[397] = 684;
        test_data[397] = 33'd7157475801;
        test_addr[398] = 199;
        test_data[398] = 33'd2378011170;
        test_addr[399] = 200;
        test_data[399] = 33'd4250933843;
        test_addr[400] = 201;
        test_data[400] = 33'd8012068873;
        test_addr[401] = 202;
        test_data[401] = 33'd2638317033;
        test_addr[402] = 203;
        test_data[402] = 33'd998547257;
        test_addr[403] = 204;
        test_data[403] = 33'd2620591812;
        test_addr[404] = 205;
        test_data[404] = 33'd2964469971;
        test_addr[405] = 113;
        test_data[405] = 33'd4144529833;
        test_addr[406] = 114;
        test_data[406] = 33'd2554819996;
        test_addr[407] = 115;
        test_data[407] = 33'd5416713673;
        test_addr[408] = 116;
        test_data[408] = 33'd1512917393;
        test_addr[409] = 117;
        test_data[409] = 33'd8261719444;
        test_addr[410] = 118;
        test_data[410] = 33'd2078089603;
        test_addr[411] = 119;
        test_data[411] = 33'd7834175968;
        test_addr[412] = 120;
        test_data[412] = 33'd5327857792;
        test_addr[413] = 121;
        test_data[413] = 33'd557179377;
        test_addr[414] = 122;
        test_data[414] = 33'd886188703;
        test_addr[415] = 123;
        test_data[415] = 33'd7600775601;
        test_addr[416] = 124;
        test_data[416] = 33'd2261534157;
        test_addr[417] = 125;
        test_data[417] = 33'd4704660590;
        test_addr[418] = 126;
        test_data[418] = 33'd717632510;
        test_addr[419] = 127;
        test_data[419] = 33'd1836818636;
        test_addr[420] = 128;
        test_data[420] = 33'd4085576191;
        test_addr[421] = 129;
        test_data[421] = 33'd5629802625;
        test_addr[422] = 130;
        test_data[422] = 33'd2760717433;
        test_addr[423] = 131;
        test_data[423] = 33'd3219734873;
        test_addr[424] = 206;
        test_data[424] = 33'd5625109385;
        test_addr[425] = 207;
        test_data[425] = 33'd155196010;
        test_addr[426] = 208;
        test_data[426] = 33'd6351840218;
        test_addr[427] = 209;
        test_data[427] = 33'd3667029732;
        test_addr[428] = 210;
        test_data[428] = 33'd7432269272;
        test_addr[429] = 211;
        test_data[429] = 33'd2875926310;
        test_addr[430] = 212;
        test_data[430] = 33'd2392747211;
        test_addr[431] = 214;
        test_data[431] = 33'd6456642822;
        test_addr[432] = 215;
        test_data[432] = 33'd8321851453;
        test_addr[433] = 216;
        test_data[433] = 33'd4576108390;
        test_addr[434] = 217;
        test_data[434] = 33'd1119239002;
        test_addr[435] = 213;
        test_data[435] = 33'd2959424098;
        test_addr[436] = 214;
        test_data[436] = 33'd2161675526;
        test_addr[437] = 215;
        test_data[437] = 33'd4026884157;
        test_addr[438] = 216;
        test_data[438] = 33'd281141094;
        test_addr[439] = 217;
        test_data[439] = 33'd1119239002;
        test_addr[440] = 218;
        test_data[440] = 33'd2296008684;
        test_addr[441] = 219;
        test_data[441] = 33'd5989901469;
        test_addr[442] = 220;
        test_data[442] = 33'd1671321966;
        test_addr[443] = 221;
        test_data[443] = 33'd1801818893;
        test_addr[444] = 222;
        test_data[444] = 33'd727510908;
        test_addr[445] = 223;
        test_data[445] = 33'd2764688405;
        test_addr[446] = 224;
        test_data[446] = 33'd2327022084;
        test_addr[447] = 225;
        test_data[447] = 33'd3019194714;
        test_addr[448] = 226;
        test_data[448] = 33'd4281849382;
        test_addr[449] = 227;
        test_data[449] = 33'd1667423717;
        test_addr[450] = 228;
        test_data[450] = 33'd4341676671;
        test_addr[451] = 229;
        test_data[451] = 33'd1506219133;
        test_addr[452] = 230;
        test_data[452] = 33'd3332009274;
        test_addr[453] = 231;
        test_data[453] = 33'd1787072800;
        test_addr[454] = 232;
        test_data[454] = 33'd6178941795;
        test_addr[455] = 233;
        test_data[455] = 33'd4512692927;
        test_addr[456] = 234;
        test_data[456] = 33'd797215018;
        test_addr[457] = 235;
        test_data[457] = 33'd3439453128;
        test_addr[458] = 236;
        test_data[458] = 33'd3012409940;
        test_addr[459] = 728;
        test_data[459] = 33'd2130178182;
        test_addr[460] = 729;
        test_data[460] = 33'd5771808161;
        test_addr[461] = 730;
        test_data[461] = 33'd3961431253;
        test_addr[462] = 731;
        test_data[462] = 33'd3189626759;
        test_addr[463] = 732;
        test_data[463] = 33'd999882873;
        test_addr[464] = 733;
        test_data[464] = 33'd5621463267;
        test_addr[465] = 734;
        test_data[465] = 33'd2715359325;
        test_addr[466] = 735;
        test_data[466] = 33'd3254548139;
        test_addr[467] = 736;
        test_data[467] = 33'd5362007932;
        test_addr[468] = 737;
        test_data[468] = 33'd2707504632;
        test_addr[469] = 738;
        test_data[469] = 33'd5608906586;
        test_addr[470] = 739;
        test_data[470] = 33'd4733897563;
        test_addr[471] = 740;
        test_data[471] = 33'd3202433012;
        test_addr[472] = 741;
        test_data[472] = 33'd6365405589;
        test_addr[473] = 742;
        test_data[473] = 33'd5582482414;
        test_addr[474] = 743;
        test_data[474] = 33'd7733373192;
        test_addr[475] = 744;
        test_data[475] = 33'd2404663132;
        test_addr[476] = 745;
        test_data[476] = 33'd4333005053;
        test_addr[477] = 746;
        test_data[477] = 33'd1546724884;
        test_addr[478] = 747;
        test_data[478] = 33'd3215049412;
        test_addr[479] = 748;
        test_data[479] = 33'd5480215175;
        test_addr[480] = 749;
        test_data[480] = 33'd6800145555;
        test_addr[481] = 750;
        test_data[481] = 33'd3873234694;
        test_addr[482] = 751;
        test_data[482] = 33'd2207759834;
        test_addr[483] = 752;
        test_data[483] = 33'd1391868779;
        test_addr[484] = 753;
        test_data[484] = 33'd5973102829;
        test_addr[485] = 754;
        test_data[485] = 33'd5229527418;
        test_addr[486] = 755;
        test_data[486] = 33'd6461474207;
        test_addr[487] = 756;
        test_data[487] = 33'd7593117400;
        test_addr[488] = 757;
        test_data[488] = 33'd2524440412;
        test_addr[489] = 758;
        test_data[489] = 33'd1681383457;
        test_addr[490] = 759;
        test_data[490] = 33'd6177082505;
        test_addr[491] = 760;
        test_data[491] = 33'd2966775552;
        test_addr[492] = 761;
        test_data[492] = 33'd6642320608;
        test_addr[493] = 762;
        test_data[493] = 33'd2301973470;
        test_addr[494] = 763;
        test_data[494] = 33'd5732931626;
        test_addr[495] = 764;
        test_data[495] = 33'd1805789468;
        test_addr[496] = 765;
        test_data[496] = 33'd1817152200;
        test_addr[497] = 766;
        test_data[497] = 33'd7417927169;
        test_addr[498] = 237;
        test_data[498] = 33'd5678123706;
        test_addr[499] = 238;
        test_data[499] = 33'd5031186309;
        test_addr[500] = 239;
        test_data[500] = 33'd3601678559;
        test_addr[501] = 240;
        test_data[501] = 33'd272401660;
        test_addr[502] = 241;
        test_data[502] = 33'd1202615656;
        test_addr[503] = 242;
        test_data[503] = 33'd7210935410;
        test_addr[504] = 243;
        test_data[504] = 33'd2004278974;
        test_addr[505] = 244;
        test_data[505] = 33'd1146573824;
        test_addr[506] = 245;
        test_data[506] = 33'd139315422;
        test_addr[507] = 246;
        test_data[507] = 33'd348319993;
        test_addr[508] = 215;
        test_data[508] = 33'd4026884157;
        test_addr[509] = 216;
        test_data[509] = 33'd6970861759;
        test_addr[510] = 247;
        test_data[510] = 33'd1238703566;
        test_addr[511] = 248;
        test_data[511] = 33'd3541486229;
        test_addr[512] = 249;
        test_data[512] = 33'd230942795;
        test_addr[513] = 250;
        test_data[513] = 33'd157822933;
        test_addr[514] = 251;
        test_data[514] = 33'd2172745435;
        test_addr[515] = 252;
        test_data[515] = 33'd3216848485;
        test_addr[516] = 253;
        test_data[516] = 33'd522192966;
        test_addr[517] = 254;
        test_data[517] = 33'd7142478840;
        test_addr[518] = 255;
        test_data[518] = 33'd714439378;
        test_addr[519] = 256;
        test_data[519] = 33'd2800244347;
        test_addr[520] = 257;
        test_data[520] = 33'd7727779294;
        test_addr[521] = 258;
        test_data[521] = 33'd3876914063;
        test_addr[522] = 259;
        test_data[522] = 33'd5457020260;
        test_addr[523] = 260;
        test_data[523] = 33'd1766135903;
        test_addr[524] = 261;
        test_data[524] = 33'd6544982435;
        test_addr[525] = 262;
        test_data[525] = 33'd5890843974;
        test_addr[526] = 263;
        test_data[526] = 33'd2114950029;
        test_addr[527] = 264;
        test_data[527] = 33'd823241581;
        test_addr[528] = 867;
        test_data[528] = 33'd11628468;
        test_addr[529] = 868;
        test_data[529] = 33'd5113552097;
        test_addr[530] = 265;
        test_data[530] = 33'd1728145956;
        test_addr[531] = 266;
        test_data[531] = 33'd6479216582;
        test_addr[532] = 267;
        test_data[532] = 33'd6336420775;
        test_addr[533] = 268;
        test_data[533] = 33'd1602773367;
        test_addr[534] = 269;
        test_data[534] = 33'd3034594309;
        test_addr[535] = 270;
        test_data[535] = 33'd5223165708;
        test_addr[536] = 271;
        test_data[536] = 33'd2102264294;
        test_addr[537] = 272;
        test_data[537] = 33'd7386511385;
        test_addr[538] = 273;
        test_data[538] = 33'd3691999146;
        test_addr[539] = 274;
        test_data[539] = 33'd2004368579;
        test_addr[540] = 275;
        test_data[540] = 33'd1824795164;
        test_addr[541] = 276;
        test_data[541] = 33'd1921721343;
        test_addr[542] = 277;
        test_data[542] = 33'd1860688658;
        test_addr[543] = 278;
        test_data[543] = 33'd7744662944;
        test_addr[544] = 279;
        test_data[544] = 33'd1883857597;
        test_addr[545] = 280;
        test_data[545] = 33'd2299961408;
        test_addr[546] = 281;
        test_data[546] = 33'd4110926899;
        test_addr[547] = 282;
        test_data[547] = 33'd8505739281;
        test_addr[548] = 283;
        test_data[548] = 33'd6894194761;
        test_addr[549] = 284;
        test_data[549] = 33'd6193308940;
        test_addr[550] = 285;
        test_data[550] = 33'd6769132966;
        test_addr[551] = 286;
        test_data[551] = 33'd775168527;
        test_addr[552] = 287;
        test_data[552] = 33'd2682374959;
        test_addr[553] = 288;
        test_data[553] = 33'd1151781196;
        test_addr[554] = 289;
        test_data[554] = 33'd6325284444;
        test_addr[555] = 290;
        test_data[555] = 33'd7978875163;
        test_addr[556] = 291;
        test_data[556] = 33'd1297973981;
        test_addr[557] = 292;
        test_data[557] = 33'd7404894283;
        test_addr[558] = 293;
        test_data[558] = 33'd688835068;
        test_addr[559] = 294;
        test_data[559] = 33'd3604100589;
        test_addr[560] = 295;
        test_data[560] = 33'd2347942712;
        test_addr[561] = 296;
        test_data[561] = 33'd1233127960;
        test_addr[562] = 297;
        test_data[562] = 33'd3955483560;
        test_addr[563] = 298;
        test_data[563] = 33'd703519346;
        test_addr[564] = 299;
        test_data[564] = 33'd8446346909;
        test_addr[565] = 300;
        test_data[565] = 33'd1320963640;
        test_addr[566] = 301;
        test_data[566] = 33'd2660948838;
        test_addr[567] = 302;
        test_data[567] = 33'd1512656212;
        test_addr[568] = 303;
        test_data[568] = 33'd7749733419;
        test_addr[569] = 304;
        test_data[569] = 33'd5311974780;
        test_addr[570] = 305;
        test_data[570] = 33'd2556845885;
        test_addr[571] = 306;
        test_data[571] = 33'd621355406;
        test_addr[572] = 307;
        test_data[572] = 33'd4594063620;
        test_addr[573] = 308;
        test_data[573] = 33'd3983220710;
        test_addr[574] = 309;
        test_data[574] = 33'd3373852337;
        test_addr[575] = 588;
        test_data[575] = 33'd1568993292;
        test_addr[576] = 589;
        test_data[576] = 33'd6590852798;
        test_addr[577] = 590;
        test_data[577] = 33'd3186803448;
        test_addr[578] = 591;
        test_data[578] = 33'd720614045;
        test_addr[579] = 592;
        test_data[579] = 33'd1698532447;
        test_addr[580] = 593;
        test_data[580] = 33'd3272624999;
        test_addr[581] = 594;
        test_data[581] = 33'd2517975264;
        test_addr[582] = 595;
        test_data[582] = 33'd6215639410;
        test_addr[583] = 310;
        test_data[583] = 33'd6937437521;
        test_addr[584] = 311;
        test_data[584] = 33'd2927272024;
        test_addr[585] = 312;
        test_data[585] = 33'd3915746261;
        test_addr[586] = 313;
        test_data[586] = 33'd494624070;
        test_addr[587] = 314;
        test_data[587] = 33'd3309988311;
        test_addr[588] = 264;
        test_data[588] = 33'd823241581;
        test_addr[589] = 265;
        test_data[589] = 33'd1728145956;
        test_addr[590] = 315;
        test_data[590] = 33'd1132837972;
        test_addr[591] = 316;
        test_data[591] = 33'd2910487772;
        test_addr[592] = 317;
        test_data[592] = 33'd4861787108;
        test_addr[593] = 318;
        test_data[593] = 33'd3655450011;
        test_addr[594] = 319;
        test_data[594] = 33'd7339518876;
        test_addr[595] = 320;
        test_data[595] = 33'd6292727298;
        test_addr[596] = 321;
        test_data[596] = 33'd7235477503;
        test_addr[597] = 322;
        test_data[597] = 33'd5267955797;
        test_addr[598] = 323;
        test_data[598] = 33'd1549846123;
        test_addr[599] = 324;
        test_data[599] = 33'd1485894970;
        test_addr[600] = 819;
        test_data[600] = 33'd3916228144;
        test_addr[601] = 820;
        test_data[601] = 33'd3676412073;
        test_addr[602] = 821;
        test_data[602] = 33'd707615435;
        test_addr[603] = 822;
        test_data[603] = 33'd661016934;
        test_addr[604] = 823;
        test_data[604] = 33'd4008531324;
        test_addr[605] = 824;
        test_data[605] = 33'd397224463;
        test_addr[606] = 825;
        test_data[606] = 33'd276834200;
        test_addr[607] = 826;
        test_data[607] = 33'd251042263;
        test_addr[608] = 827;
        test_data[608] = 33'd8085273827;
        test_addr[609] = 828;
        test_data[609] = 33'd3353314327;
        test_addr[610] = 829;
        test_data[610] = 33'd4734411430;
        test_addr[611] = 325;
        test_data[611] = 33'd1503820403;
        test_addr[612] = 326;
        test_data[612] = 33'd20706691;
        test_addr[613] = 327;
        test_data[613] = 33'd8038799687;
        test_addr[614] = 328;
        test_data[614] = 33'd5940114068;
        test_addr[615] = 329;
        test_data[615] = 33'd6225941925;
        test_addr[616] = 330;
        test_data[616] = 33'd1408921763;
        test_addr[617] = 343;
        test_data[617] = 33'd7509816123;
        test_addr[618] = 344;
        test_data[618] = 33'd3796226835;
        test_addr[619] = 345;
        test_data[619] = 33'd3794021488;
        test_addr[620] = 346;
        test_data[620] = 33'd7472813135;
        test_addr[621] = 347;
        test_data[621] = 33'd5644318223;
        test_addr[622] = 348;
        test_data[622] = 33'd5382171239;
        test_addr[623] = 349;
        test_data[623] = 33'd7979830920;
        test_addr[624] = 350;
        test_data[624] = 33'd1629934311;
        test_addr[625] = 351;
        test_data[625] = 33'd3124014635;
        test_addr[626] = 352;
        test_data[626] = 33'd3793842303;
        test_addr[627] = 353;
        test_data[627] = 33'd5449735842;
        test_addr[628] = 354;
        test_data[628] = 33'd701425537;
        test_addr[629] = 355;
        test_data[629] = 33'd5673958092;
        test_addr[630] = 356;
        test_data[630] = 33'd2020066253;
        test_addr[631] = 357;
        test_data[631] = 33'd2661076722;
        test_addr[632] = 358;
        test_data[632] = 33'd2161533557;
        test_addr[633] = 359;
        test_data[633] = 33'd2495672481;
        test_addr[634] = 360;
        test_data[634] = 33'd1452465810;
        test_addr[635] = 331;
        test_data[635] = 33'd1012710083;
        test_addr[636] = 332;
        test_data[636] = 33'd3964024451;
        test_addr[637] = 333;
        test_data[637] = 33'd5314426613;
        test_addr[638] = 334;
        test_data[638] = 33'd1631873129;
        test_addr[639] = 335;
        test_data[639] = 33'd3094982513;
        test_addr[640] = 336;
        test_data[640] = 33'd604229382;
        test_addr[641] = 337;
        test_data[641] = 33'd190701906;
        test_addr[642] = 338;
        test_data[642] = 33'd2063414812;
        test_addr[643] = 339;
        test_data[643] = 33'd2384267827;
        test_addr[644] = 340;
        test_data[644] = 33'd2877406934;
        test_addr[645] = 341;
        test_data[645] = 33'd2186863965;
        test_addr[646] = 342;
        test_data[646] = 33'd4078357046;
        test_addr[647] = 343;
        test_data[647] = 33'd3214848827;
        test_addr[648] = 344;
        test_data[648] = 33'd3796226835;
        test_addr[649] = 345;
        test_data[649] = 33'd5984959799;
        test_addr[650] = 346;
        test_data[650] = 33'd3177845839;
        test_addr[651] = 347;
        test_data[651] = 33'd1349350927;
        test_addr[652] = 348;
        test_data[652] = 33'd6200100403;
        test_addr[653] = 1;
        test_data[653] = 33'd1897396466;
        test_addr[654] = 2;
        test_data[654] = 33'd1865453439;
        test_addr[655] = 3;
        test_data[655] = 33'd1011693257;
        test_addr[656] = 4;
        test_data[656] = 33'd93557296;
        test_addr[657] = 5;
        test_data[657] = 33'd838687445;
        test_addr[658] = 6;
        test_data[658] = 33'd3274300910;
        test_addr[659] = 7;
        test_data[659] = 33'd3491080214;
        test_addr[660] = 8;
        test_data[660] = 33'd5725858811;
        test_addr[661] = 349;
        test_data[661] = 33'd3684863624;
        test_addr[662] = 350;
        test_data[662] = 33'd1629934311;
        test_addr[663] = 351;
        test_data[663] = 33'd3124014635;
        test_addr[664] = 352;
        test_data[664] = 33'd7842412105;
        test_addr[665] = 353;
        test_data[665] = 33'd7669866197;
        test_addr[666] = 354;
        test_data[666] = 33'd701425537;
        test_addr[667] = 355;
        test_data[667] = 33'd1378990796;
        test_addr[668] = 356;
        test_data[668] = 33'd2020066253;
        test_addr[669] = 440;
        test_data[669] = 33'd5225182815;
        test_addr[670] = 441;
        test_data[670] = 33'd4133778867;
        test_addr[671] = 442;
        test_data[671] = 33'd1182124915;
        test_addr[672] = 443;
        test_data[672] = 33'd887054320;
        test_addr[673] = 444;
        test_data[673] = 33'd3362594900;
        test_addr[674] = 445;
        test_data[674] = 33'd6136562966;
        test_addr[675] = 446;
        test_data[675] = 33'd2862511605;
        test_addr[676] = 447;
        test_data[676] = 33'd2384680284;
        test_addr[677] = 448;
        test_data[677] = 33'd1262035775;
        test_addr[678] = 449;
        test_data[678] = 33'd8095724258;
        test_addr[679] = 357;
        test_data[679] = 33'd7527261121;
        test_addr[680] = 358;
        test_data[680] = 33'd2161533557;
        test_addr[681] = 359;
        test_data[681] = 33'd2495672481;
        test_addr[682] = 161;
        test_data[682] = 33'd3824367798;
        test_addr[683] = 162;
        test_data[683] = 33'd1461900145;
        test_addr[684] = 163;
        test_data[684] = 33'd2334826380;
        test_addr[685] = 164;
        test_data[685] = 33'd617221806;
        test_addr[686] = 165;
        test_data[686] = 33'd117310100;
        test_addr[687] = 166;
        test_data[687] = 33'd2648221725;
        test_addr[688] = 360;
        test_data[688] = 33'd1452465810;
        test_addr[689] = 361;
        test_data[689] = 33'd3160518389;
        test_addr[690] = 362;
        test_data[690] = 33'd2841382309;
        test_addr[691] = 363;
        test_data[691] = 33'd6519326376;
        test_addr[692] = 364;
        test_data[692] = 33'd2996693876;
        test_addr[693] = 509;
        test_data[693] = 33'd2012699169;
        test_addr[694] = 510;
        test_data[694] = 33'd8373460279;
        test_addr[695] = 511;
        test_data[695] = 33'd868517225;
        test_addr[696] = 512;
        test_data[696] = 33'd3892061908;
        test_addr[697] = 365;
        test_data[697] = 33'd4840238116;
        test_addr[698] = 366;
        test_data[698] = 33'd3707227066;
        test_addr[699] = 367;
        test_data[699] = 33'd1471019555;
        test_addr[700] = 479;
        test_data[700] = 33'd3609861208;
        test_addr[701] = 480;
        test_data[701] = 33'd1712226038;
        test_addr[702] = 481;
        test_data[702] = 33'd6192543376;
        test_addr[703] = 482;
        test_data[703] = 33'd3069633443;
        test_addr[704] = 483;
        test_data[704] = 33'd2649187208;
        test_addr[705] = 484;
        test_data[705] = 33'd4269737784;
        test_addr[706] = 485;
        test_data[706] = 33'd3345226134;
        test_addr[707] = 486;
        test_data[707] = 33'd5619184823;
        test_addr[708] = 487;
        test_data[708] = 33'd4754141521;
        test_addr[709] = 488;
        test_data[709] = 33'd7405527561;
        test_addr[710] = 489;
        test_data[710] = 33'd1491360199;
        test_addr[711] = 490;
        test_data[711] = 33'd1608490784;
        test_addr[712] = 491;
        test_data[712] = 33'd1594847873;
        test_addr[713] = 492;
        test_data[713] = 33'd5581589871;
        test_addr[714] = 493;
        test_data[714] = 33'd1800880124;
        test_addr[715] = 494;
        test_data[715] = 33'd821347042;
        test_addr[716] = 368;
        test_data[716] = 33'd5865918636;
        test_addr[717] = 369;
        test_data[717] = 33'd2915294719;
        test_addr[718] = 370;
        test_data[718] = 33'd1041307001;
        test_addr[719] = 371;
        test_data[719] = 33'd2929810272;
        test_addr[720] = 372;
        test_data[720] = 33'd6496116180;
        test_addr[721] = 373;
        test_data[721] = 33'd5625508504;
        test_addr[722] = 374;
        test_data[722] = 33'd86209782;
        test_addr[723] = 375;
        test_data[723] = 33'd6196947805;
        test_addr[724] = 376;
        test_data[724] = 33'd2739596899;
        test_addr[725] = 377;
        test_data[725] = 33'd528252277;
        test_addr[726] = 378;
        test_data[726] = 33'd1303994115;
        test_addr[727] = 571;
        test_data[727] = 33'd2590447935;
        test_addr[728] = 572;
        test_data[728] = 33'd8195598141;
        test_addr[729] = 573;
        test_data[729] = 33'd4029761842;
        test_addr[730] = 574;
        test_data[730] = 33'd4104262188;
        test_addr[731] = 575;
        test_data[731] = 33'd197152237;
        test_addr[732] = 576;
        test_data[732] = 33'd65320894;
        test_addr[733] = 577;
        test_data[733] = 33'd4153629096;
        test_addr[734] = 578;
        test_data[734] = 33'd741309116;
        test_addr[735] = 579;
        test_data[735] = 33'd8196884014;
        test_addr[736] = 580;
        test_data[736] = 33'd3021320586;
        test_addr[737] = 379;
        test_data[737] = 33'd7784253901;
        test_addr[738] = 380;
        test_data[738] = 33'd909919624;
        test_addr[739] = 857;
        test_data[739] = 33'd2231454879;
        test_addr[740] = 858;
        test_data[740] = 33'd4000613725;
        test_addr[741] = 859;
        test_data[741] = 33'd544317971;
        test_addr[742] = 860;
        test_data[742] = 33'd7040706922;
        test_addr[743] = 861;
        test_data[743] = 33'd1495467381;
        test_addr[744] = 862;
        test_data[744] = 33'd3532219985;
        test_addr[745] = 381;
        test_data[745] = 33'd2494821825;
        test_addr[746] = 382;
        test_data[746] = 33'd2070296687;
        test_addr[747] = 383;
        test_data[747] = 33'd489544890;
        test_addr[748] = 384;
        test_data[748] = 33'd6082388754;
        test_addr[749] = 385;
        test_data[749] = 33'd8460081423;
        test_addr[750] = 386;
        test_data[750] = 33'd1757687415;
        test_addr[751] = 387;
        test_data[751] = 33'd3967144044;
        test_addr[752] = 388;
        test_data[752] = 33'd2794749959;
        test_addr[753] = 389;
        test_data[753] = 33'd3611635867;
        test_addr[754] = 390;
        test_data[754] = 33'd1980103462;
        test_addr[755] = 391;
        test_data[755] = 33'd7007931198;
        test_addr[756] = 392;
        test_data[756] = 33'd1088256129;
        test_addr[757] = 393;
        test_data[757] = 33'd2750675278;
        test_addr[758] = 394;
        test_data[758] = 33'd862789604;
        test_addr[759] = 395;
        test_data[759] = 33'd2126893221;
        test_addr[760] = 396;
        test_data[760] = 33'd4286897536;
        test_addr[761] = 397;
        test_data[761] = 33'd1575257700;
        test_addr[762] = 476;
        test_data[762] = 33'd3314836530;
        test_addr[763] = 477;
        test_data[763] = 33'd2300423720;
        test_addr[764] = 478;
        test_data[764] = 33'd3938658140;
        test_addr[765] = 479;
        test_data[765] = 33'd3609861208;
        test_addr[766] = 480;
        test_data[766] = 33'd1712226038;
        test_addr[767] = 481;
        test_data[767] = 33'd1897576080;
        test_addr[768] = 482;
        test_data[768] = 33'd3069633443;
        test_addr[769] = 483;
        test_data[769] = 33'd2649187208;
        test_addr[770] = 484;
        test_data[770] = 33'd4269737784;
        test_addr[771] = 398;
        test_data[771] = 33'd3564413496;
        test_addr[772] = 399;
        test_data[772] = 33'd8348795707;
        test_addr[773] = 400;
        test_data[773] = 33'd523664291;
        test_addr[774] = 401;
        test_data[774] = 33'd6146695502;
        test_addr[775] = 402;
        test_data[775] = 33'd7337650168;
        test_addr[776] = 403;
        test_data[776] = 33'd3751867044;
        test_addr[777] = 404;
        test_data[777] = 33'd478746838;
        test_addr[778] = 405;
        test_data[778] = 33'd5510167281;
        test_addr[779] = 406;
        test_data[779] = 33'd272467445;
        test_addr[780] = 407;
        test_data[780] = 33'd7206734832;
        test_addr[781] = 408;
        test_data[781] = 33'd4272217241;
        test_addr[782] = 409;
        test_data[782] = 33'd2962982112;
        test_addr[783] = 435;
        test_data[783] = 33'd4337287957;
        test_addr[784] = 436;
        test_data[784] = 33'd3478059314;
        test_addr[785] = 437;
        test_data[785] = 33'd6918768709;
        test_addr[786] = 438;
        test_data[786] = 33'd5301336794;
        test_addr[787] = 439;
        test_data[787] = 33'd4263494862;
        test_addr[788] = 440;
        test_data[788] = 33'd930215519;
        test_addr[789] = 441;
        test_data[789] = 33'd4133778867;
        test_addr[790] = 442;
        test_data[790] = 33'd1182124915;
        test_addr[791] = 443;
        test_data[791] = 33'd4974900993;
        test_addr[792] = 444;
        test_data[792] = 33'd3362594900;
        test_addr[793] = 445;
        test_data[793] = 33'd8315861511;
        test_addr[794] = 446;
        test_data[794] = 33'd2862511605;
        test_addr[795] = 447;
        test_data[795] = 33'd6891560402;
        test_addr[796] = 448;
        test_data[796] = 33'd5288579862;
        test_addr[797] = 449;
        test_data[797] = 33'd3800756962;
        test_addr[798] = 450;
        test_data[798] = 33'd3977574422;
        test_addr[799] = 451;
        test_data[799] = 33'd3943760075;
        test_addr[800] = 452;
        test_data[800] = 33'd4807830;
        test_addr[801] = 453;
        test_data[801] = 33'd6015439001;
        test_addr[802] = 454;
        test_data[802] = 33'd2119829098;
        test_addr[803] = 455;
        test_data[803] = 33'd6260016904;
        test_addr[804] = 456;
        test_data[804] = 33'd2711175043;
        test_addr[805] = 457;
        test_data[805] = 33'd2493892019;
        test_addr[806] = 458;
        test_data[806] = 33'd5198951104;
        test_addr[807] = 459;
        test_data[807] = 33'd600779198;
        test_addr[808] = 460;
        test_data[808] = 33'd2977339794;
        test_addr[809] = 461;
        test_data[809] = 33'd4758217052;
        test_addr[810] = 410;
        test_data[810] = 33'd327705331;
        test_addr[811] = 411;
        test_data[811] = 33'd1638656261;
        test_addr[812] = 90;
        test_data[812] = 33'd7824485414;
        test_addr[813] = 91;
        test_data[813] = 33'd1285586415;
        test_addr[814] = 92;
        test_data[814] = 33'd2746581280;
        test_addr[815] = 93;
        test_data[815] = 33'd3760806334;
        test_addr[816] = 94;
        test_data[816] = 33'd2987649344;
        test_addr[817] = 95;
        test_data[817] = 33'd2737991781;
        test_addr[818] = 96;
        test_data[818] = 33'd7927622917;
        test_addr[819] = 412;
        test_data[819] = 33'd1831501086;
        test_addr[820] = 413;
        test_data[820] = 33'd3893899942;
        test_addr[821] = 414;
        test_data[821] = 33'd1927908942;
        test_addr[822] = 415;
        test_data[822] = 33'd3159116717;
        test_addr[823] = 416;
        test_data[823] = 33'd5514170026;
        test_addr[824] = 417;
        test_data[824] = 33'd2072738163;
        test_addr[825] = 418;
        test_data[825] = 33'd717648603;
        test_addr[826] = 419;
        test_data[826] = 33'd2628348997;
        test_addr[827] = 420;
        test_data[827] = 33'd8205518102;
        test_addr[828] = 421;
        test_data[828] = 33'd1376576240;
        test_addr[829] = 422;
        test_data[829] = 33'd712524200;
        test_addr[830] = 423;
        test_data[830] = 33'd3658904312;
        test_addr[831] = 424;
        test_data[831] = 33'd6352407140;
        test_addr[832] = 425;
        test_data[832] = 33'd4239458745;
        test_addr[833] = 426;
        test_data[833] = 33'd5813495832;
        test_addr[834] = 427;
        test_data[834] = 33'd6612773170;
        test_addr[835] = 428;
        test_data[835] = 33'd3161887892;
        test_addr[836] = 429;
        test_data[836] = 33'd523036013;
        test_addr[837] = 430;
        test_data[837] = 33'd4102642570;
        test_addr[838] = 431;
        test_data[838] = 33'd4615300648;
        test_addr[839] = 432;
        test_data[839] = 33'd1817537658;
        test_addr[840] = 433;
        test_data[840] = 33'd131728541;
        test_addr[841] = 434;
        test_data[841] = 33'd4343734793;
        test_addr[842] = 435;
        test_data[842] = 33'd8148602079;
        test_addr[843] = 436;
        test_data[843] = 33'd3478059314;
        test_addr[844] = 437;
        test_data[844] = 33'd2623801413;
        test_addr[845] = 438;
        test_data[845] = 33'd1006369498;
        test_addr[846] = 439;
        test_data[846] = 33'd4263494862;
        test_addr[847] = 440;
        test_data[847] = 33'd5126970118;
        test_addr[848] = 441;
        test_data[848] = 33'd4339589118;
        test_addr[849] = 442;
        test_data[849] = 33'd1182124915;
        test_addr[850] = 443;
        test_data[850] = 33'd7399585677;
        test_addr[851] = 444;
        test_data[851] = 33'd6385755315;
        test_addr[852] = 445;
        test_data[852] = 33'd4020894215;
        test_addr[853] = 446;
        test_data[853] = 33'd2862511605;
        test_addr[854] = 447;
        test_data[854] = 33'd7605716756;
        test_addr[855] = 448;
        test_data[855] = 33'd8042654791;
        test_addr[856] = 449;
        test_data[856] = 33'd3800756962;
        test_addr[857] = 450;
        test_data[857] = 33'd3977574422;
        test_addr[858] = 451;
        test_data[858] = 33'd3943760075;
        test_addr[859] = 452;
        test_data[859] = 33'd4638952883;
        test_addr[860] = 453;
        test_data[860] = 33'd1720471705;
        test_addr[861] = 454;
        test_data[861] = 33'd7595125484;
        test_addr[862] = 455;
        test_data[862] = 33'd5690363224;
        test_addr[863] = 456;
        test_data[863] = 33'd2711175043;
        test_addr[864] = 457;
        test_data[864] = 33'd2493892019;
        test_addr[865] = 458;
        test_data[865] = 33'd903983808;
        test_addr[866] = 459;
        test_data[866] = 33'd600779198;
        test_addr[867] = 460;
        test_data[867] = 33'd6932226628;
        test_addr[868] = 461;
        test_data[868] = 33'd463249756;
        test_addr[869] = 462;
        test_data[869] = 33'd1387176348;
        test_addr[870] = 463;
        test_data[870] = 33'd4096796069;
        test_addr[871] = 464;
        test_data[871] = 33'd1087715771;
        test_addr[872] = 465;
        test_data[872] = 33'd2637855582;
        test_addr[873] = 466;
        test_data[873] = 33'd2023239053;
        test_addr[874] = 467;
        test_data[874] = 33'd579888698;
        test_addr[875] = 468;
        test_data[875] = 33'd4524566999;
        test_addr[876] = 469;
        test_data[876] = 33'd3850513177;
        test_addr[877] = 470;
        test_data[877] = 33'd8053591198;
        test_addr[878] = 471;
        test_data[878] = 33'd8572755322;
        test_addr[879] = 472;
        test_data[879] = 33'd5391691702;
        test_addr[880] = 473;
        test_data[880] = 33'd7236249197;
        test_addr[881] = 474;
        test_data[881] = 33'd4051137299;
        test_addr[882] = 228;
        test_data[882] = 33'd46709375;
        test_addr[883] = 229;
        test_data[883] = 33'd1506219133;
        test_addr[884] = 230;
        test_data[884] = 33'd3332009274;
        test_addr[885] = 231;
        test_data[885] = 33'd1787072800;
        test_addr[886] = 232;
        test_data[886] = 33'd1883974499;
        test_addr[887] = 233;
        test_data[887] = 33'd7252466501;
        test_addr[888] = 475;
        test_data[888] = 33'd3259448472;
        test_addr[889] = 476;
        test_data[889] = 33'd3314836530;
        test_addr[890] = 477;
        test_data[890] = 33'd2300423720;
        test_addr[891] = 478;
        test_data[891] = 33'd3938658140;
        test_addr[892] = 479;
        test_data[892] = 33'd5700204836;
        test_addr[893] = 480;
        test_data[893] = 33'd1712226038;
        test_addr[894] = 481;
        test_data[894] = 33'd8251203677;
        test_addr[895] = 482;
        test_data[895] = 33'd3069633443;
        test_addr[896] = 483;
        test_data[896] = 33'd2649187208;
        test_addr[897] = 484;
        test_data[897] = 33'd4269737784;
        test_addr[898] = 485;
        test_data[898] = 33'd3345226134;
        test_addr[899] = 486;
        test_data[899] = 33'd1324217527;
        test_addr[900] = 487;
        test_data[900] = 33'd459174225;
        test_addr[901] = 488;
        test_data[901] = 33'd4766687662;
        test_addr[902] = 489;
        test_data[902] = 33'd1491360199;
        test_addr[903] = 490;
        test_data[903] = 33'd7509750402;
        test_addr[904] = 491;
        test_data[904] = 33'd7840319602;
        test_addr[905] = 492;
        test_data[905] = 33'd5140269978;
        test_addr[906] = 493;
        test_data[906] = 33'd1800880124;
        test_addr[907] = 494;
        test_data[907] = 33'd821347042;
        test_addr[908] = 495;
        test_data[908] = 33'd2117462048;
        test_addr[909] = 496;
        test_data[909] = 33'd3581785694;
        test_addr[910] = 497;
        test_data[910] = 33'd1177368502;
        test_addr[911] = 498;
        test_data[911] = 33'd3822144455;
        test_addr[912] = 499;
        test_data[912] = 33'd3127083966;
        test_addr[913] = 63;
        test_data[913] = 33'd6375058737;
        test_addr[914] = 64;
        test_data[914] = 33'd4280548596;
        test_addr[915] = 65;
        test_data[915] = 33'd3000665519;
        test_addr[916] = 66;
        test_data[916] = 33'd2358437066;
        test_addr[917] = 67;
        test_data[917] = 33'd1974385293;
        test_addr[918] = 68;
        test_data[918] = 33'd4811908333;
        test_addr[919] = 69;
        test_data[919] = 33'd6399762141;
        test_addr[920] = 70;
        test_data[920] = 33'd8002874760;
        test_addr[921] = 500;
        test_data[921] = 33'd6256130330;
        test_addr[922] = 501;
        test_data[922] = 33'd4890683210;
        test_addr[923] = 502;
        test_data[923] = 33'd1457378795;
        test_addr[924] = 503;
        test_data[924] = 33'd3251093126;
        test_addr[925] = 504;
        test_data[925] = 33'd2586581290;
        test_addr[926] = 505;
        test_data[926] = 33'd2328699311;
        test_addr[927] = 506;
        test_data[927] = 33'd6484913381;
        test_addr[928] = 507;
        test_data[928] = 33'd5085193235;
        test_addr[929] = 508;
        test_data[929] = 33'd5045897300;
        test_addr[930] = 509;
        test_data[930] = 33'd4867108699;
        test_addr[931] = 510;
        test_data[931] = 33'd6033729221;
        test_addr[932] = 511;
        test_data[932] = 33'd868517225;
        test_addr[933] = 512;
        test_data[933] = 33'd7929692789;
        test_addr[934] = 513;
        test_data[934] = 33'd45075662;
        test_addr[935] = 514;
        test_data[935] = 33'd3808305303;
        test_addr[936] = 515;
        test_data[936] = 33'd934899158;
        test_addr[937] = 516;
        test_data[937] = 33'd7572361486;
        test_addr[938] = 914;
        test_data[938] = 33'd617611722;
        test_addr[939] = 915;
        test_data[939] = 33'd316048180;
        test_addr[940] = 916;
        test_data[940] = 33'd5255126288;
        test_addr[941] = 917;
        test_data[941] = 33'd347883434;
        test_addr[942] = 918;
        test_data[942] = 33'd1901704297;
        test_addr[943] = 919;
        test_data[943] = 33'd1993211956;
        test_addr[944] = 920;
        test_data[944] = 33'd1049468648;
        test_addr[945] = 921;
        test_data[945] = 33'd4539358254;
        test_addr[946] = 922;
        test_data[946] = 33'd268862713;
        test_addr[947] = 923;
        test_data[947] = 33'd2554414221;
        test_addr[948] = 924;
        test_data[948] = 33'd5459260817;
        test_addr[949] = 925;
        test_data[949] = 33'd74622926;
        test_addr[950] = 926;
        test_data[950] = 33'd2262293352;
        test_addr[951] = 927;
        test_data[951] = 33'd4526097193;
        test_addr[952] = 517;
        test_data[952] = 33'd5559008313;
        test_addr[953] = 518;
        test_data[953] = 33'd209533787;
        test_addr[954] = 519;
        test_data[954] = 33'd2029500360;
        test_addr[955] = 520;
        test_data[955] = 33'd6245576239;
        test_addr[956] = 521;
        test_data[956] = 33'd5463034538;
        test_addr[957] = 522;
        test_data[957] = 33'd6324429409;
        test_addr[958] = 523;
        test_data[958] = 33'd3215894844;
        test_addr[959] = 524;
        test_data[959] = 33'd8015135462;
        test_addr[960] = 525;
        test_data[960] = 33'd2968836141;
        test_addr[961] = 526;
        test_data[961] = 33'd2513327218;
        test_addr[962] = 527;
        test_data[962] = 33'd3681101907;
        test_addr[963] = 79;
        test_data[963] = 33'd4395530772;
        test_addr[964] = 528;
        test_data[964] = 33'd1983832739;
        test_addr[965] = 529;
        test_data[965] = 33'd3177420342;
        test_addr[966] = 530;
        test_data[966] = 33'd4972277676;
        test_addr[967] = 576;
        test_data[967] = 33'd65320894;
        test_addr[968] = 577;
        test_data[968] = 33'd4153629096;
        test_addr[969] = 578;
        test_data[969] = 33'd741309116;
        test_addr[970] = 579;
        test_data[970] = 33'd7581792795;
        test_addr[971] = 580;
        test_data[971] = 33'd5978452235;
        test_addr[972] = 581;
        test_data[972] = 33'd2322605034;
        test_addr[973] = 582;
        test_data[973] = 33'd3186320755;
        test_addr[974] = 583;
        test_data[974] = 33'd2141613643;
        test_addr[975] = 531;
        test_data[975] = 33'd4269338406;
        test_addr[976] = 532;
        test_data[976] = 33'd1758387349;
        test_addr[977] = 533;
        test_data[977] = 33'd3892039782;
        test_addr[978] = 534;
        test_data[978] = 33'd8425250671;
        test_addr[979] = 535;
        test_data[979] = 33'd335471988;
        test_addr[980] = 536;
        test_data[980] = 33'd3377477922;
        test_addr[981] = 537;
        test_data[981] = 33'd6752854290;
        test_addr[982] = 538;
        test_data[982] = 33'd1250172866;
        test_addr[983] = 539;
        test_data[983] = 33'd7821327008;
        test_addr[984] = 540;
        test_data[984] = 33'd7780906832;
        test_addr[985] = 541;
        test_data[985] = 33'd8338169444;
        test_addr[986] = 542;
        test_data[986] = 33'd7570455396;
        test_addr[987] = 543;
        test_data[987] = 33'd6343418035;
        test_addr[988] = 544;
        test_data[988] = 33'd2034855529;
        test_addr[989] = 545;
        test_data[989] = 33'd4717977195;
        test_addr[990] = 546;
        test_data[990] = 33'd5361340914;
        test_addr[991] = 547;
        test_data[991] = 33'd3961698218;
        test_addr[992] = 548;
        test_data[992] = 33'd3807612461;
        test_addr[993] = 549;
        test_data[993] = 33'd2484022925;
        test_addr[994] = 550;
        test_data[994] = 33'd2131016181;
        test_addr[995] = 551;
        test_data[995] = 33'd4294945315;
        test_addr[996] = 552;
        test_data[996] = 33'd3583226745;
        test_addr[997] = 553;
        test_data[997] = 33'd81343249;
        test_addr[998] = 554;
        test_data[998] = 33'd7619314565;
        test_addr[999] = 555;
        test_data[999] = 33'd3198658539;
        test_addr[1000] = 257;
        test_data[1000] = 33'd7372178857;
        test_addr[1001] = 258;
        test_data[1001] = 33'd3876914063;
        test_addr[1002] = 259;
        test_data[1002] = 33'd5086348149;
        test_addr[1003] = 260;
        test_data[1003] = 33'd1766135903;
        test_addr[1004] = 261;
        test_data[1004] = 33'd2250015139;
        test_addr[1005] = 262;
        test_data[1005] = 33'd8041716152;
        test_addr[1006] = 263;
        test_data[1006] = 33'd2114950029;
        test_addr[1007] = 264;
        test_data[1007] = 33'd6030676047;
        test_addr[1008] = 265;
        test_data[1008] = 33'd1728145956;
        test_addr[1009] = 266;
        test_data[1009] = 33'd5475497812;
        test_addr[1010] = 556;
        test_data[1010] = 33'd174607435;
        test_addr[1011] = 557;
        test_data[1011] = 33'd1596273533;
        test_addr[1012] = 558;
        test_data[1012] = 33'd862985215;
        test_addr[1013] = 559;
        test_data[1013] = 33'd7206462729;
        test_addr[1014] = 560;
        test_data[1014] = 33'd4558624291;
        test_addr[1015] = 561;
        test_data[1015] = 33'd2008701872;
        test_addr[1016] = 562;
        test_data[1016] = 33'd1056483800;
        test_addr[1017] = 563;
        test_data[1017] = 33'd5765863846;
        test_addr[1018] = 564;
        test_data[1018] = 33'd5005038697;
        test_addr[1019] = 565;
        test_data[1019] = 33'd8319482882;
        test_addr[1020] = 566;
        test_data[1020] = 33'd1836238996;
        test_addr[1021] = 567;
        test_data[1021] = 33'd5187007025;
        test_addr[1022] = 568;
        test_data[1022] = 33'd2411940668;
        test_addr[1023] = 38;
        test_data[1023] = 33'd4595738108;
        test_addr[1024] = 39;
        test_data[1024] = 33'd1715945728;
        test_addr[1025] = 569;
        test_data[1025] = 33'd2786633091;
        test_addr[1026] = 537;
        test_data[1026] = 33'd2457886994;
        test_addr[1027] = 538;
        test_data[1027] = 33'd1250172866;
        test_addr[1028] = 539;
        test_data[1028] = 33'd3526359712;
        test_addr[1029] = 540;
        test_data[1029] = 33'd3485939536;
        test_addr[1030] = 541;
        test_data[1030] = 33'd7130223703;
        test_addr[1031] = 542;
        test_data[1031] = 33'd7918912706;
        test_addr[1032] = 570;
        test_data[1032] = 33'd5028079524;
        test_addr[1033] = 571;
        test_data[1033] = 33'd2590447935;
        test_addr[1034] = 572;
        test_data[1034] = 33'd3900630845;
        test_addr[1035] = 573;
        test_data[1035] = 33'd6062395255;
        test_addr[1036] = 574;
        test_data[1036] = 33'd4104262188;
        test_addr[1037] = 575;
        test_data[1037] = 33'd197152237;
        test_addr[1038] = 576;
        test_data[1038] = 33'd65320894;
        test_addr[1039] = 654;
        test_data[1039] = 33'd1955032163;
        test_addr[1040] = 655;
        test_data[1040] = 33'd3509997369;
        test_addr[1041] = 656;
        test_data[1041] = 33'd5144493049;
        test_addr[1042] = 657;
        test_data[1042] = 33'd4073638024;
        test_addr[1043] = 658;
        test_data[1043] = 33'd420911824;
        test_addr[1044] = 659;
        test_data[1044] = 33'd5214547350;
        test_addr[1045] = 660;
        test_data[1045] = 33'd270341019;
        test_addr[1046] = 577;
        test_data[1046] = 33'd7487456487;
        test_addr[1047] = 303;
        test_data[1047] = 33'd3454766123;
        test_addr[1048] = 304;
        test_data[1048] = 33'd1017007484;
        test_addr[1049] = 305;
        test_data[1049] = 33'd2556845885;
        test_addr[1050] = 306;
        test_data[1050] = 33'd621355406;
        test_addr[1051] = 307;
        test_data[1051] = 33'd299096324;
        test_addr[1052] = 308;
        test_data[1052] = 33'd3983220710;
        test_addr[1053] = 309;
        test_data[1053] = 33'd3373852337;
        test_addr[1054] = 310;
        test_data[1054] = 33'd8366721803;
        test_addr[1055] = 311;
        test_data[1055] = 33'd7453268996;
        test_addr[1056] = 312;
        test_data[1056] = 33'd3915746261;
        test_addr[1057] = 313;
        test_data[1057] = 33'd494624070;
        test_addr[1058] = 314;
        test_data[1058] = 33'd3309988311;
        test_addr[1059] = 315;
        test_data[1059] = 33'd1132837972;
        test_addr[1060] = 316;
        test_data[1060] = 33'd7155650735;
        test_addr[1061] = 317;
        test_data[1061] = 33'd566819812;
        test_addr[1062] = 318;
        test_data[1062] = 33'd3655450011;
        test_addr[1063] = 319;
        test_data[1063] = 33'd3044551580;
        test_addr[1064] = 320;
        test_data[1064] = 33'd1997760002;
        test_addr[1065] = 321;
        test_data[1065] = 33'd2940510207;
        test_addr[1066] = 322;
        test_data[1066] = 33'd6770792044;
        test_addr[1067] = 323;
        test_data[1067] = 33'd1549846123;
        test_addr[1068] = 578;
        test_data[1068] = 33'd741309116;
        test_addr[1069] = 579;
        test_data[1069] = 33'd3286825499;
        test_addr[1070] = 580;
        test_data[1070] = 33'd4437226894;
        test_addr[1071] = 581;
        test_data[1071] = 33'd6786210540;
        test_addr[1072] = 582;
        test_data[1072] = 33'd3186320755;
        test_addr[1073] = 583;
        test_data[1073] = 33'd5546564331;
        test_addr[1074] = 584;
        test_data[1074] = 33'd7021976841;
        test_addr[1075] = 585;
        test_data[1075] = 33'd1415357636;
        test_addr[1076] = 586;
        test_data[1076] = 33'd3407577517;
        test_addr[1077] = 587;
        test_data[1077] = 33'd976124543;
        test_addr[1078] = 588;
        test_data[1078] = 33'd1568993292;
        test_addr[1079] = 589;
        test_data[1079] = 33'd2295885502;
        test_addr[1080] = 590;
        test_data[1080] = 33'd4965483023;
        test_addr[1081] = 591;
        test_data[1081] = 33'd720614045;
        test_addr[1082] = 592;
        test_data[1082] = 33'd4962358397;
        test_addr[1083] = 593;
        test_data[1083] = 33'd3272624999;
        test_addr[1084] = 594;
        test_data[1084] = 33'd6298732118;
        test_addr[1085] = 595;
        test_data[1085] = 33'd1920672114;
        test_addr[1086] = 596;
        test_data[1086] = 33'd5712487399;
        test_addr[1087] = 597;
        test_data[1087] = 33'd2479920114;
        test_addr[1088] = 598;
        test_data[1088] = 33'd4421365779;
        test_addr[1089] = 599;
        test_data[1089] = 33'd8047374456;
        test_addr[1090] = 600;
        test_data[1090] = 33'd3556822102;
        test_addr[1091] = 601;
        test_data[1091] = 33'd750890938;
        test_addr[1092] = 273;
        test_data[1092] = 33'd3691999146;
        test_addr[1093] = 274;
        test_data[1093] = 33'd5110340957;
        test_addr[1094] = 275;
        test_data[1094] = 33'd1824795164;
        test_addr[1095] = 276;
        test_data[1095] = 33'd7954072775;
        test_addr[1096] = 277;
        test_data[1096] = 33'd7836451389;
        test_addr[1097] = 278;
        test_data[1097] = 33'd6725185953;
        test_addr[1098] = 279;
        test_data[1098] = 33'd1883857597;
        test_addr[1099] = 280;
        test_data[1099] = 33'd8133671110;
        test_addr[1100] = 281;
        test_data[1100] = 33'd4864858501;
        test_addr[1101] = 282;
        test_data[1101] = 33'd7125549996;
        test_addr[1102] = 283;
        test_data[1102] = 33'd7399715496;
        test_addr[1103] = 284;
        test_data[1103] = 33'd7700695726;
        test_addr[1104] = 285;
        test_data[1104] = 33'd2474165670;
        test_addr[1105] = 286;
        test_data[1105] = 33'd775168527;
        test_addr[1106] = 287;
        test_data[1106] = 33'd2682374959;
        test_addr[1107] = 288;
        test_data[1107] = 33'd1151781196;
        test_addr[1108] = 289;
        test_data[1108] = 33'd2030317148;
        test_addr[1109] = 290;
        test_data[1109] = 33'd8539951632;
        test_addr[1110] = 291;
        test_data[1110] = 33'd1297973981;
        test_addr[1111] = 292;
        test_data[1111] = 33'd3109926987;
        test_addr[1112] = 602;
        test_data[1112] = 33'd5291659124;
        test_addr[1113] = 603;
        test_data[1113] = 33'd7333581249;
        test_addr[1114] = 604;
        test_data[1114] = 33'd8402652528;
        test_addr[1115] = 605;
        test_data[1115] = 33'd4062492645;
        test_addr[1116] = 606;
        test_data[1116] = 33'd3682415596;
        test_addr[1117] = 607;
        test_data[1117] = 33'd7003166823;
        test_addr[1118] = 608;
        test_data[1118] = 33'd4965065868;
        test_addr[1119] = 609;
        test_data[1119] = 33'd412456713;
        test_addr[1120] = 610;
        test_data[1120] = 33'd3240265434;
        test_addr[1121] = 611;
        test_data[1121] = 33'd3431050438;
        test_addr[1122] = 612;
        test_data[1122] = 33'd551188312;
        test_addr[1123] = 613;
        test_data[1123] = 33'd3036714220;
        test_addr[1124] = 614;
        test_data[1124] = 33'd1362451819;
        test_addr[1125] = 615;
        test_data[1125] = 33'd3586907395;
        test_addr[1126] = 616;
        test_data[1126] = 33'd1633853584;
        test_addr[1127] = 617;
        test_data[1127] = 33'd404883268;
        test_addr[1128] = 618;
        test_data[1128] = 33'd7131734700;
        test_addr[1129] = 619;
        test_data[1129] = 33'd3850720077;
        test_addr[1130] = 620;
        test_data[1130] = 33'd6863363118;
        test_addr[1131] = 621;
        test_data[1131] = 33'd5954122527;
        test_addr[1132] = 265;
        test_data[1132] = 33'd1728145956;
        test_addr[1133] = 266;
        test_data[1133] = 33'd4762901115;
        test_addr[1134] = 267;
        test_data[1134] = 33'd2041453479;
        test_addr[1135] = 268;
        test_data[1135] = 33'd1602773367;
        test_addr[1136] = 269;
        test_data[1136] = 33'd3034594309;
        test_addr[1137] = 270;
        test_data[1137] = 33'd7801331469;
        test_addr[1138] = 271;
        test_data[1138] = 33'd2102264294;
        test_addr[1139] = 272;
        test_data[1139] = 33'd7282734714;
        test_addr[1140] = 273;
        test_data[1140] = 33'd3691999146;
        test_addr[1141] = 274;
        test_data[1141] = 33'd4814273926;
        test_addr[1142] = 275;
        test_data[1142] = 33'd4411654374;
        test_addr[1143] = 276;
        test_data[1143] = 33'd5502431853;
        test_addr[1144] = 277;
        test_data[1144] = 33'd6996885009;
        test_addr[1145] = 278;
        test_data[1145] = 33'd2430218657;
        test_addr[1146] = 279;
        test_data[1146] = 33'd5475402475;
        test_addr[1147] = 280;
        test_data[1147] = 33'd7017824608;
        test_addr[1148] = 281;
        test_data[1148] = 33'd569891205;
        test_addr[1149] = 282;
        test_data[1149] = 33'd6634607199;
        test_addr[1150] = 283;
        test_data[1150] = 33'd3104748200;
        test_addr[1151] = 284;
        test_data[1151] = 33'd3405728430;
        test_addr[1152] = 285;
        test_data[1152] = 33'd2474165670;
        test_addr[1153] = 286;
        test_data[1153] = 33'd775168527;
        test_addr[1154] = 287;
        test_data[1154] = 33'd2682374959;
        test_addr[1155] = 288;
        test_data[1155] = 33'd1151781196;
        test_addr[1156] = 289;
        test_data[1156] = 33'd6696644380;
        test_addr[1157] = 622;
        test_data[1157] = 33'd5233181935;
        test_addr[1158] = 623;
        test_data[1158] = 33'd1096932212;
        test_addr[1159] = 624;
        test_data[1159] = 33'd1317201626;
        test_addr[1160] = 625;
        test_data[1160] = 33'd1251593008;
        test_addr[1161] = 626;
        test_data[1161] = 33'd3713789991;
        test_addr[1162] = 627;
        test_data[1162] = 33'd1679511367;
        test_addr[1163] = 628;
        test_data[1163] = 33'd3449788833;
        test_addr[1164] = 629;
        test_data[1164] = 33'd1317727169;
        test_addr[1165] = 630;
        test_data[1165] = 33'd3548473177;
        test_addr[1166] = 631;
        test_data[1166] = 33'd2390103675;
        test_addr[1167] = 632;
        test_data[1167] = 33'd173501673;
        test_addr[1168] = 633;
        test_data[1168] = 33'd2419434228;
        test_addr[1169] = 634;
        test_data[1169] = 33'd6846033658;
        test_addr[1170] = 635;
        test_data[1170] = 33'd8061767602;
        test_addr[1171] = 636;
        test_data[1171] = 33'd130031873;
        test_addr[1172] = 637;
        test_data[1172] = 33'd7231712843;
        test_addr[1173] = 848;
        test_data[1173] = 33'd1989148088;
        test_addr[1174] = 849;
        test_data[1174] = 33'd4029825875;
        test_addr[1175] = 850;
        test_data[1175] = 33'd3859470178;
        test_addr[1176] = 851;
        test_data[1176] = 33'd3497740514;
        test_addr[1177] = 638;
        test_data[1177] = 33'd8497020465;
        test_addr[1178] = 66;
        test_data[1178] = 33'd2358437066;
        test_addr[1179] = 67;
        test_data[1179] = 33'd1974385293;
        test_addr[1180] = 68;
        test_data[1180] = 33'd516941037;
        test_addr[1181] = 69;
        test_data[1181] = 33'd6229536401;
        test_addr[1182] = 70;
        test_data[1182] = 33'd5045883796;
        test_addr[1183] = 71;
        test_data[1183] = 33'd2915912397;
        test_addr[1184] = 72;
        test_data[1184] = 33'd1456092511;
        test_addr[1185] = 73;
        test_data[1185] = 33'd3301388465;
        test_addr[1186] = 74;
        test_data[1186] = 33'd8247363629;
        test_addr[1187] = 75;
        test_data[1187] = 33'd2806077644;
        test_addr[1188] = 76;
        test_data[1188] = 33'd2442953578;
        test_addr[1189] = 77;
        test_data[1189] = 33'd2962067559;
        test_addr[1190] = 78;
        test_data[1190] = 33'd2225443136;
        test_addr[1191] = 79;
        test_data[1191] = 33'd100563476;
        test_addr[1192] = 80;
        test_data[1192] = 33'd3727744700;
        test_addr[1193] = 81;
        test_data[1193] = 33'd7123838722;
        test_addr[1194] = 82;
        test_data[1194] = 33'd1564001926;
        test_addr[1195] = 639;
        test_data[1195] = 33'd2378925636;
        test_addr[1196] = 640;
        test_data[1196] = 33'd2328757272;
        test_addr[1197] = 641;
        test_data[1197] = 33'd6543107895;
        test_addr[1198] = 642;
        test_data[1198] = 33'd8466757322;
        test_addr[1199] = 643;
        test_data[1199] = 33'd5193322176;
        test_addr[1200] = 644;
        test_data[1200] = 33'd487448243;
        test_addr[1201] = 645;
        test_data[1201] = 33'd1218724220;
        test_addr[1202] = 646;
        test_data[1202] = 33'd1152709717;
        test_addr[1203] = 734;
        test_data[1203] = 33'd5577659723;
        test_addr[1204] = 735;
        test_data[1204] = 33'd3254548139;
        test_addr[1205] = 736;
        test_data[1205] = 33'd5033134688;
        test_addr[1206] = 737;
        test_data[1206] = 33'd6690819010;
        test_addr[1207] = 738;
        test_data[1207] = 33'd1313939290;
        test_addr[1208] = 739;
        test_data[1208] = 33'd438930267;
        test_addr[1209] = 740;
        test_data[1209] = 33'd3202433012;
        test_addr[1210] = 741;
        test_data[1210] = 33'd5246498121;
        test_addr[1211] = 742;
        test_data[1211] = 33'd4644948962;
        test_addr[1212] = 743;
        test_data[1212] = 33'd7382275344;
        test_addr[1213] = 744;
        test_data[1213] = 33'd2404663132;
        test_addr[1214] = 745;
        test_data[1214] = 33'd4297256878;
        test_addr[1215] = 746;
        test_data[1215] = 33'd1546724884;
        test_addr[1216] = 747;
        test_data[1216] = 33'd3215049412;
        test_addr[1217] = 748;
        test_data[1217] = 33'd1185247879;
        test_addr[1218] = 749;
        test_data[1218] = 33'd2505178259;
        test_addr[1219] = 750;
        test_data[1219] = 33'd3873234694;
        test_addr[1220] = 751;
        test_data[1220] = 33'd2207759834;
        test_addr[1221] = 752;
        test_data[1221] = 33'd1391868779;
        test_addr[1222] = 753;
        test_data[1222] = 33'd1678135533;
        test_addr[1223] = 754;
        test_data[1223] = 33'd934560122;
        test_addr[1224] = 755;
        test_data[1224] = 33'd2166506911;
        test_addr[1225] = 756;
        test_data[1225] = 33'd3298150104;
        test_addr[1226] = 647;
        test_data[1226] = 33'd6422156778;
        test_addr[1227] = 648;
        test_data[1227] = 33'd776883759;
        test_addr[1228] = 649;
        test_data[1228] = 33'd3154846827;
        test_addr[1229] = 650;
        test_data[1229] = 33'd1968337716;
        test_addr[1230] = 651;
        test_data[1230] = 33'd2766237222;
        test_addr[1231] = 652;
        test_data[1231] = 33'd1737322648;
        test_addr[1232] = 653;
        test_data[1232] = 33'd3358716186;
        test_addr[1233] = 654;
        test_data[1233] = 33'd1955032163;
        test_addr[1234] = 655;
        test_data[1234] = 33'd3509997369;
        test_addr[1235] = 656;
        test_data[1235] = 33'd5198895715;
        test_addr[1236] = 657;
        test_data[1236] = 33'd4073638024;
        test_addr[1237] = 658;
        test_data[1237] = 33'd420911824;
        test_addr[1238] = 659;
        test_data[1238] = 33'd4826581421;
        test_addr[1239] = 660;
        test_data[1239] = 33'd5996206537;
        test_addr[1240] = 661;
        test_data[1240] = 33'd3720845072;
        test_addr[1241] = 662;
        test_data[1241] = 33'd2741441705;
        test_addr[1242] = 663;
        test_data[1242] = 33'd4758750375;
        test_addr[1243] = 664;
        test_data[1243] = 33'd961409848;
        test_addr[1244] = 665;
        test_data[1244] = 33'd3437855889;
        test_addr[1245] = 666;
        test_data[1245] = 33'd3656350260;
        test_addr[1246] = 667;
        test_data[1246] = 33'd8039394718;
        test_addr[1247] = 668;
        test_data[1247] = 33'd2346181448;
        test_addr[1248] = 669;
        test_data[1248] = 33'd8162854371;
        test_addr[1249] = 670;
        test_data[1249] = 33'd4565285525;
        test_addr[1250] = 671;
        test_data[1250] = 33'd660543359;
        test_addr[1251] = 672;
        test_data[1251] = 33'd3657343727;
        test_addr[1252] = 673;
        test_data[1252] = 33'd8380808575;
        test_addr[1253] = 674;
        test_data[1253] = 33'd1495437377;
        test_addr[1254] = 675;
        test_data[1254] = 33'd3828766155;
        test_addr[1255] = 676;
        test_data[1255] = 33'd1442188537;
        test_addr[1256] = 677;
        test_data[1256] = 33'd4176733826;
        test_addr[1257] = 678;
        test_data[1257] = 33'd2975839092;
        test_addr[1258] = 679;
        test_data[1258] = 33'd1411385993;
        test_addr[1259] = 680;
        test_data[1259] = 33'd4893901514;
        test_addr[1260] = 681;
        test_data[1260] = 33'd3370337054;
        test_addr[1261] = 682;
        test_data[1261] = 33'd180214976;
        test_addr[1262] = 683;
        test_data[1262] = 33'd452619150;
        test_addr[1263] = 684;
        test_data[1263] = 33'd2862508505;
        test_addr[1264] = 685;
        test_data[1264] = 33'd4501609240;
        test_addr[1265] = 797;
        test_data[1265] = 33'd3852826982;
        test_addr[1266] = 798;
        test_data[1266] = 33'd1995026993;
        test_addr[1267] = 799;
        test_data[1267] = 33'd3803697363;
        test_addr[1268] = 800;
        test_data[1268] = 33'd3694851582;
        test_addr[1269] = 686;
        test_data[1269] = 33'd3310495543;
        test_addr[1270] = 687;
        test_data[1270] = 33'd7386678733;
        test_addr[1271] = 673;
        test_data[1271] = 33'd4085841279;
        test_addr[1272] = 674;
        test_data[1272] = 33'd1495437377;
        test_addr[1273] = 675;
        test_data[1273] = 33'd3828766155;
        test_addr[1274] = 676;
        test_data[1274] = 33'd4831963502;
        test_addr[1275] = 677;
        test_data[1275] = 33'd4176733826;
        test_addr[1276] = 678;
        test_data[1276] = 33'd2975839092;
        test_addr[1277] = 679;
        test_data[1277] = 33'd4914535390;
        test_addr[1278] = 680;
        test_data[1278] = 33'd598934218;
        test_addr[1279] = 681;
        test_data[1279] = 33'd3370337054;
        test_addr[1280] = 682;
        test_data[1280] = 33'd180214976;
        test_addr[1281] = 683;
        test_data[1281] = 33'd452619150;
        test_addr[1282] = 688;
        test_data[1282] = 33'd3075220499;
        test_addr[1283] = 689;
        test_data[1283] = 33'd1724620145;
        test_addr[1284] = 690;
        test_data[1284] = 33'd3106437015;
        test_addr[1285] = 691;
        test_data[1285] = 33'd3982442458;
        test_addr[1286] = 692;
        test_data[1286] = 33'd1622816285;
        test_addr[1287] = 693;
        test_data[1287] = 33'd3113725398;
        test_addr[1288] = 694;
        test_data[1288] = 33'd62309893;
        test_addr[1289] = 155;
        test_data[1289] = 33'd3182442945;
        test_addr[1290] = 156;
        test_data[1290] = 33'd4176867573;
        test_addr[1291] = 157;
        test_data[1291] = 33'd6881806575;
        test_addr[1292] = 158;
        test_data[1292] = 33'd6193217737;
        test_addr[1293] = 159;
        test_data[1293] = 33'd2928595937;
        test_addr[1294] = 160;
        test_data[1294] = 33'd660917259;
        test_addr[1295] = 161;
        test_data[1295] = 33'd4818269575;
        test_addr[1296] = 162;
        test_data[1296] = 33'd1461900145;
        test_addr[1297] = 163;
        test_data[1297] = 33'd2334826380;
        test_addr[1298] = 164;
        test_data[1298] = 33'd8537771313;
        test_addr[1299] = 165;
        test_data[1299] = 33'd117310100;
        test_addr[1300] = 166;
        test_data[1300] = 33'd4583374828;
        test_addr[1301] = 167;
        test_data[1301] = 33'd3641515376;
        test_addr[1302] = 168;
        test_data[1302] = 33'd5817113770;
        test_addr[1303] = 169;
        test_data[1303] = 33'd4949526821;
        test_addr[1304] = 695;
        test_data[1304] = 33'd7208943391;
        test_addr[1305] = 696;
        test_data[1305] = 33'd274861910;
        test_addr[1306] = 697;
        test_data[1306] = 33'd3794458561;
        test_addr[1307] = 698;
        test_data[1307] = 33'd154010637;
        test_addr[1308] = 699;
        test_data[1308] = 33'd3680508728;
        test_addr[1309] = 700;
        test_data[1309] = 33'd1353090612;
        test_addr[1310] = 701;
        test_data[1310] = 33'd3933897631;
        test_addr[1311] = 702;
        test_data[1311] = 33'd1901550375;
        test_addr[1312] = 703;
        test_data[1312] = 33'd2171400527;
        test_addr[1313] = 704;
        test_data[1313] = 33'd5308682605;
        test_addr[1314] = 705;
        test_data[1314] = 33'd1050986732;
        test_addr[1315] = 706;
        test_data[1315] = 33'd8018341824;
        test_addr[1316] = 707;
        test_data[1316] = 33'd2518819451;
        test_addr[1317] = 708;
        test_data[1317] = 33'd3912899891;
        test_addr[1318] = 709;
        test_data[1318] = 33'd8165083887;
        test_addr[1319] = 710;
        test_data[1319] = 33'd5575708910;
        test_addr[1320] = 711;
        test_data[1320] = 33'd2022344989;
        test_addr[1321] = 712;
        test_data[1321] = 33'd1962337977;
        test_addr[1322] = 713;
        test_data[1322] = 33'd3785505943;
        test_addr[1323] = 714;
        test_data[1323] = 33'd7705198144;
        test_addr[1324] = 715;
        test_data[1324] = 33'd8264211677;
        test_addr[1325] = 716;
        test_data[1325] = 33'd1756901617;
        test_addr[1326] = 717;
        test_data[1326] = 33'd6957447495;
        test_addr[1327] = 718;
        test_data[1327] = 33'd4730160309;
        test_addr[1328] = 719;
        test_data[1328] = 33'd7580694984;
        test_addr[1329] = 720;
        test_data[1329] = 33'd6521262767;
        test_addr[1330] = 721;
        test_data[1330] = 33'd3305804503;
        test_addr[1331] = 722;
        test_data[1331] = 33'd3177944058;
        test_addr[1332] = 723;
        test_data[1332] = 33'd1900853036;
        test_addr[1333] = 724;
        test_data[1333] = 33'd3326485598;
        test_addr[1334] = 725;
        test_data[1334] = 33'd1069406399;
        test_addr[1335] = 726;
        test_data[1335] = 33'd4007895896;
        test_addr[1336] = 727;
        test_data[1336] = 33'd2861577116;
        test_addr[1337] = 728;
        test_data[1337] = 33'd2130178182;
        test_addr[1338] = 729;
        test_data[1338] = 33'd1476840865;
        test_addr[1339] = 730;
        test_data[1339] = 33'd3961431253;
        test_addr[1340] = 731;
        test_data[1340] = 33'd5611763044;
        test_addr[1341] = 732;
        test_data[1341] = 33'd4409825708;
        test_addr[1342] = 733;
        test_data[1342] = 33'd5592431471;
        test_addr[1343] = 910;
        test_data[1343] = 33'd5420224974;
        test_addr[1344] = 911;
        test_data[1344] = 33'd7934725460;
        test_addr[1345] = 912;
        test_data[1345] = 33'd1323603140;
        test_addr[1346] = 734;
        test_data[1346] = 33'd1282692427;
        test_addr[1347] = 735;
        test_data[1347] = 33'd3254548139;
        test_addr[1348] = 736;
        test_data[1348] = 33'd738167392;
        test_addr[1349] = 737;
        test_data[1349] = 33'd8376832557;
        test_addr[1350] = 738;
        test_data[1350] = 33'd1313939290;
        test_addr[1351] = 430;
        test_data[1351] = 33'd4102642570;
        test_addr[1352] = 431;
        test_data[1352] = 33'd4540922993;
        test_addr[1353] = 432;
        test_data[1353] = 33'd1817537658;
        test_addr[1354] = 433;
        test_data[1354] = 33'd131728541;
        test_addr[1355] = 434;
        test_data[1355] = 33'd48767497;
        test_addr[1356] = 435;
        test_data[1356] = 33'd4366891633;
        test_addr[1357] = 436;
        test_data[1357] = 33'd3478059314;
        test_addr[1358] = 437;
        test_data[1358] = 33'd2623801413;
        test_addr[1359] = 438;
        test_data[1359] = 33'd7022976476;
        test_addr[1360] = 739;
        test_data[1360] = 33'd438930267;
        test_addr[1361] = 740;
        test_data[1361] = 33'd3202433012;
        test_addr[1362] = 741;
        test_data[1362] = 33'd951530825;
        test_addr[1363] = 742;
        test_data[1363] = 33'd349981666;
        test_addr[1364] = 890;
        test_data[1364] = 33'd1018830267;
        test_addr[1365] = 891;
        test_data[1365] = 33'd4197184161;
        test_addr[1366] = 892;
        test_data[1366] = 33'd1771063249;
        test_addr[1367] = 893;
        test_data[1367] = 33'd2729806528;
        test_addr[1368] = 894;
        test_data[1368] = 33'd1657957379;
        test_addr[1369] = 895;
        test_data[1369] = 33'd1344756801;
        test_addr[1370] = 743;
        test_data[1370] = 33'd3087308048;
        test_addr[1371] = 744;
        test_data[1371] = 33'd2404663132;
        test_addr[1372] = 745;
        test_data[1372] = 33'd2289582;
        test_addr[1373] = 746;
        test_data[1373] = 33'd1546724884;
        test_addr[1374] = 747;
        test_data[1374] = 33'd3215049412;
        test_addr[1375] = 748;
        test_data[1375] = 33'd1185247879;
        test_addr[1376] = 749;
        test_data[1376] = 33'd2505178259;
        test_addr[1377] = 750;
        test_data[1377] = 33'd8024259215;
        test_addr[1378] = 751;
        test_data[1378] = 33'd5599021950;
        test_addr[1379] = 752;
        test_data[1379] = 33'd1391868779;
        test_addr[1380] = 753;
        test_data[1380] = 33'd1678135533;
        test_addr[1381] = 754;
        test_data[1381] = 33'd8469280287;
        test_addr[1382] = 755;
        test_data[1382] = 33'd2166506911;
        test_addr[1383] = 756;
        test_data[1383] = 33'd3298150104;
        test_addr[1384] = 949;
        test_data[1384] = 33'd318477808;
        test_addr[1385] = 950;
        test_data[1385] = 33'd5506740052;
        test_addr[1386] = 757;
        test_data[1386] = 33'd2524440412;
        test_addr[1387] = 758;
        test_data[1387] = 33'd5007970228;
        test_addr[1388] = 759;
        test_data[1388] = 33'd1882115209;
        test_addr[1389] = 760;
        test_data[1389] = 33'd2966775552;
        test_addr[1390] = 761;
        test_data[1390] = 33'd2347353312;
        test_addr[1391] = 762;
        test_data[1391] = 33'd2301973470;
        test_addr[1392] = 763;
        test_data[1392] = 33'd1437964330;
        test_addr[1393] = 764;
        test_data[1393] = 33'd5730676846;
        test_addr[1394] = 765;
        test_data[1394] = 33'd1817152200;
        test_addr[1395] = 766;
        test_data[1395] = 33'd3122959873;
        test_addr[1396] = 767;
        test_data[1396] = 33'd2928940173;
        test_addr[1397] = 768;
        test_data[1397] = 33'd2226595292;
        test_addr[1398] = 769;
        test_data[1398] = 33'd4489833474;
        test_addr[1399] = 770;
        test_data[1399] = 33'd968883625;
        test_addr[1400] = 771;
        test_data[1400] = 33'd1262750963;
        test_addr[1401] = 772;
        test_data[1401] = 33'd4061278725;
        test_addr[1402] = 773;
        test_data[1402] = 33'd7931842053;
        test_addr[1403] = 774;
        test_data[1403] = 33'd877880049;
        test_addr[1404] = 775;
        test_data[1404] = 33'd3939170061;
        test_addr[1405] = 776;
        test_data[1405] = 33'd2515051088;
        test_addr[1406] = 777;
        test_data[1406] = 33'd3175216081;
        test_addr[1407] = 778;
        test_data[1407] = 33'd6703764433;
        test_addr[1408] = 779;
        test_data[1408] = 33'd7514416922;
        test_addr[1409] = 780;
        test_data[1409] = 33'd2476818174;
        test_addr[1410] = 781;
        test_data[1410] = 33'd2253784569;
        test_addr[1411] = 782;
        test_data[1411] = 33'd357526767;
        test_addr[1412] = 783;
        test_data[1412] = 33'd6946993805;
        test_addr[1413] = 784;
        test_data[1413] = 33'd560379488;
        test_addr[1414] = 785;
        test_data[1414] = 33'd2691045821;
        test_addr[1415] = 786;
        test_data[1415] = 33'd8197121458;
        test_addr[1416] = 787;
        test_data[1416] = 33'd109264237;
        test_addr[1417] = 788;
        test_data[1417] = 33'd1639691474;
        test_addr[1418] = 789;
        test_data[1418] = 33'd2090407313;
        test_addr[1419] = 790;
        test_data[1419] = 33'd8271843708;
        test_addr[1420] = 791;
        test_data[1420] = 33'd496190147;
        test_addr[1421] = 792;
        test_data[1421] = 33'd8285308490;
        test_addr[1422] = 793;
        test_data[1422] = 33'd1132372465;
        test_addr[1423] = 794;
        test_data[1423] = 33'd2371798522;
        test_addr[1424] = 603;
        test_data[1424] = 33'd3038613953;
        test_addr[1425] = 604;
        test_data[1425] = 33'd5244145147;
        test_addr[1426] = 605;
        test_data[1426] = 33'd4062492645;
        test_addr[1427] = 606;
        test_data[1427] = 33'd3682415596;
        test_addr[1428] = 795;
        test_data[1428] = 33'd2253800365;
        test_addr[1429] = 796;
        test_data[1429] = 33'd1668815192;
        test_addr[1430] = 797;
        test_data[1430] = 33'd3852826982;
        test_addr[1431] = 798;
        test_data[1431] = 33'd1995026993;
        test_addr[1432] = 799;
        test_data[1432] = 33'd6918212362;
        test_addr[1433] = 800;
        test_data[1433] = 33'd3694851582;
        test_addr[1434] = 801;
        test_data[1434] = 33'd4632347571;
        test_addr[1435] = 802;
        test_data[1435] = 33'd3175044348;
        test_addr[1436] = 803;
        test_data[1436] = 33'd5314478180;
        test_addr[1437] = 804;
        test_data[1437] = 33'd8045352922;
        test_addr[1438] = 805;
        test_data[1438] = 33'd627959300;
        test_addr[1439] = 806;
        test_data[1439] = 33'd3113296974;
        test_addr[1440] = 110;
        test_data[1440] = 33'd4027024129;
        test_addr[1441] = 111;
        test_data[1441] = 33'd645329535;
        test_addr[1442] = 807;
        test_data[1442] = 33'd1709814211;
        test_addr[1443] = 808;
        test_data[1443] = 33'd3076343433;
        test_addr[1444] = 809;
        test_data[1444] = 33'd1538329166;
        test_addr[1445] = 810;
        test_data[1445] = 33'd914364136;
        test_addr[1446] = 811;
        test_data[1446] = 33'd5625369704;
        test_addr[1447] = 812;
        test_data[1447] = 33'd2940558418;
        test_addr[1448] = 813;
        test_data[1448] = 33'd5947736261;
        test_addr[1449] = 814;
        test_data[1449] = 33'd5679802670;
        test_addr[1450] = 815;
        test_data[1450] = 33'd6655695583;
        test_addr[1451] = 816;
        test_data[1451] = 33'd96275483;
        test_addr[1452] = 817;
        test_data[1452] = 33'd1666061305;
        test_addr[1453] = 818;
        test_data[1453] = 33'd160882647;
        test_addr[1454] = 819;
        test_data[1454] = 33'd3916228144;
        test_addr[1455] = 820;
        test_data[1455] = 33'd3676412073;
        test_addr[1456] = 734;
        test_data[1456] = 33'd6277313401;
        test_addr[1457] = 735;
        test_data[1457] = 33'd3254548139;
        test_addr[1458] = 736;
        test_data[1458] = 33'd738167392;
        test_addr[1459] = 821;
        test_data[1459] = 33'd707615435;
        test_addr[1460] = 271;
        test_data[1460] = 33'd2102264294;
        test_addr[1461] = 272;
        test_data[1461] = 33'd2987767418;
        test_addr[1462] = 273;
        test_data[1462] = 33'd6614304677;
        test_addr[1463] = 274;
        test_data[1463] = 33'd5964409563;
        test_addr[1464] = 275;
        test_data[1464] = 33'd5405099483;
        test_addr[1465] = 276;
        test_data[1465] = 33'd1207464557;
        test_addr[1466] = 822;
        test_data[1466] = 33'd4730189416;
        test_addr[1467] = 823;
        test_data[1467] = 33'd4008531324;
        test_addr[1468] = 824;
        test_data[1468] = 33'd5782203292;
        test_addr[1469] = 825;
        test_data[1469] = 33'd276834200;
        test_addr[1470] = 826;
        test_data[1470] = 33'd251042263;
        test_addr[1471] = 827;
        test_data[1471] = 33'd3790306531;
        test_addr[1472] = 251;
        test_data[1472] = 33'd2172745435;
        test_addr[1473] = 252;
        test_data[1473] = 33'd3216848485;
        test_addr[1474] = 253;
        test_data[1474] = 33'd522192966;
        test_addr[1475] = 254;
        test_data[1475] = 33'd2847511544;
        test_addr[1476] = 255;
        test_data[1476] = 33'd5244171905;
        test_addr[1477] = 256;
        test_data[1477] = 33'd2800244347;
        test_addr[1478] = 828;
        test_data[1478] = 33'd3353314327;
        test_addr[1479] = 829;
        test_data[1479] = 33'd6096115965;
        test_addr[1480] = 830;
        test_data[1480] = 33'd7224575749;
        test_addr[1481] = 831;
        test_data[1481] = 33'd11545355;
        test_addr[1482] = 832;
        test_data[1482] = 33'd2809961330;
        test_addr[1483] = 833;
        test_data[1483] = 33'd1455017460;
        test_addr[1484] = 834;
        test_data[1484] = 33'd6276411338;
        test_addr[1485] = 835;
        test_data[1485] = 33'd5210735480;
        test_addr[1486] = 836;
        test_data[1486] = 33'd2037704408;
        test_addr[1487] = 837;
        test_data[1487] = 33'd1657911559;
        test_addr[1488] = 838;
        test_data[1488] = 33'd924586107;
        test_addr[1489] = 839;
        test_data[1489] = 33'd1862425237;
        test_addr[1490] = 275;
        test_data[1490] = 33'd7708246555;
        test_addr[1491] = 276;
        test_data[1491] = 33'd5750505125;
        test_addr[1492] = 277;
        test_data[1492] = 33'd2701917713;
        test_addr[1493] = 278;
        test_data[1493] = 33'd2430218657;
        test_addr[1494] = 279;
        test_data[1494] = 33'd1180435179;
        test_addr[1495] = 280;
        test_data[1495] = 33'd7179835914;
        test_addr[1496] = 281;
        test_data[1496] = 33'd569891205;
        test_addr[1497] = 282;
        test_data[1497] = 33'd2339639903;
        test_addr[1498] = 283;
        test_data[1498] = 33'd4412201310;
        test_addr[1499] = 284;
        test_data[1499] = 33'd3405728430;
        test_addr[1500] = 285;
        test_data[1500] = 33'd2474165670;
        test_addr[1501] = 286;
        test_data[1501] = 33'd775168527;
        test_addr[1502] = 287;
        test_data[1502] = 33'd5726672532;
        test_addr[1503] = 288;
        test_data[1503] = 33'd1151781196;
        test_addr[1504] = 840;
        test_data[1504] = 33'd5262935972;
        test_addr[1505] = 841;
        test_data[1505] = 33'd209372675;
        test_addr[1506] = 842;
        test_data[1506] = 33'd7547394232;
        test_addr[1507] = 843;
        test_data[1507] = 33'd4105319985;
        test_addr[1508] = 844;
        test_data[1508] = 33'd4108930760;
        test_addr[1509] = 845;
        test_data[1509] = 33'd3010963361;
        test_addr[1510] = 846;
        test_data[1510] = 33'd5710490928;
        test_addr[1511] = 847;
        test_data[1511] = 33'd2811533726;
        test_addr[1512] = 848;
        test_data[1512] = 33'd1989148088;
        test_addr[1513] = 849;
        test_data[1513] = 33'd7038811373;
        test_addr[1514] = 850;
        test_data[1514] = 33'd3859470178;
        test_addr[1515] = 851;
        test_data[1515] = 33'd5831938632;
        test_addr[1516] = 852;
        test_data[1516] = 33'd7676369681;
        test_addr[1517] = 853;
        test_data[1517] = 33'd2928255153;
        test_addr[1518] = 854;
        test_data[1518] = 33'd4252373770;
        test_addr[1519] = 855;
        test_data[1519] = 33'd7943658595;
        test_addr[1520] = 856;
        test_data[1520] = 33'd3274644583;
        test_addr[1521] = 857;
        test_data[1521] = 33'd6512958584;
        test_addr[1522] = 344;
        test_data[1522] = 33'd3796226835;
        test_addr[1523] = 345;
        test_data[1523] = 33'd1689992503;
        test_addr[1524] = 858;
        test_data[1524] = 33'd4000613725;
        test_addr[1525] = 859;
        test_data[1525] = 33'd544317971;
        test_addr[1526] = 860;
        test_data[1526] = 33'd2745739626;
        test_addr[1527] = 861;
        test_data[1527] = 33'd1495467381;
        test_addr[1528] = 862;
        test_data[1528] = 33'd3532219985;
        test_addr[1529] = 863;
        test_data[1529] = 33'd6628643768;
        test_addr[1530] = 864;
        test_data[1530] = 33'd4724362607;
        test_addr[1531] = 865;
        test_data[1531] = 33'd8235096157;
        test_addr[1532] = 866;
        test_data[1532] = 33'd284044551;
        test_addr[1533] = 867;
        test_data[1533] = 33'd11628468;
        test_addr[1534] = 868;
        test_data[1534] = 33'd818584801;
        test_addr[1535] = 869;
        test_data[1535] = 33'd2050504608;
        test_addr[1536] = 870;
        test_data[1536] = 33'd2235229089;
        test_addr[1537] = 871;
        test_data[1537] = 33'd4323262799;
        test_addr[1538] = 872;
        test_data[1538] = 33'd3498935539;
        test_addr[1539] = 873;
        test_data[1539] = 33'd2783581831;
        test_addr[1540] = 874;
        test_data[1540] = 33'd3793369460;
        test_addr[1541] = 290;
        test_data[1541] = 33'd5262524120;
        test_addr[1542] = 291;
        test_data[1542] = 33'd7412524491;
        test_addr[1543] = 292;
        test_data[1543] = 33'd5721523613;
        test_addr[1544] = 293;
        test_data[1544] = 33'd688835068;
        test_addr[1545] = 294;
        test_data[1545] = 33'd4502455750;
        test_addr[1546] = 295;
        test_data[1546] = 33'd2347942712;
        test_addr[1547] = 296;
        test_data[1547] = 33'd1233127960;
        test_addr[1548] = 875;
        test_data[1548] = 33'd4043269648;
        test_addr[1549] = 876;
        test_data[1549] = 33'd1362121102;
        test_addr[1550] = 877;
        test_data[1550] = 33'd5891494679;
        test_addr[1551] = 731;
        test_data[1551] = 33'd1316795748;
        test_addr[1552] = 732;
        test_data[1552] = 33'd114858412;
        test_addr[1553] = 733;
        test_data[1553] = 33'd1297464175;
        test_addr[1554] = 734;
        test_data[1554] = 33'd1982346105;
        test_addr[1555] = 735;
        test_data[1555] = 33'd5715371284;
        test_addr[1556] = 736;
        test_data[1556] = 33'd4883711229;
        test_addr[1557] = 737;
        test_data[1557] = 33'd4081865261;
        test_addr[1558] = 738;
        test_data[1558] = 33'd1313939290;
        test_addr[1559] = 739;
        test_data[1559] = 33'd7986992125;
        test_addr[1560] = 740;
        test_data[1560] = 33'd3202433012;
        test_addr[1561] = 741;
        test_data[1561] = 33'd951530825;
        test_addr[1562] = 742;
        test_data[1562] = 33'd4902879794;
        test_addr[1563] = 743;
        test_data[1563] = 33'd3087308048;
        test_addr[1564] = 744;
        test_data[1564] = 33'd2404663132;
        test_addr[1565] = 745;
        test_data[1565] = 33'd6982470618;
        test_addr[1566] = 746;
        test_data[1566] = 33'd1546724884;
        test_addr[1567] = 747;
        test_data[1567] = 33'd5556930029;
        test_addr[1568] = 748;
        test_data[1568] = 33'd1185247879;
        test_addr[1569] = 749;
        test_data[1569] = 33'd4676430554;
        test_addr[1570] = 750;
        test_data[1570] = 33'd3729291919;
        test_addr[1571] = 751;
        test_data[1571] = 33'd1304054654;
        test_addr[1572] = 878;
        test_data[1572] = 33'd886953612;
        test_addr[1573] = 879;
        test_data[1573] = 33'd8384258756;
        test_addr[1574] = 880;
        test_data[1574] = 33'd1513837228;
        test_addr[1575] = 881;
        test_data[1575] = 33'd1205481735;
        test_addr[1576] = 882;
        test_data[1576] = 33'd6699088219;
        test_addr[1577] = 883;
        test_data[1577] = 33'd6790344467;
        test_addr[1578] = 884;
        test_data[1578] = 33'd1603698784;
        test_addr[1579] = 885;
        test_data[1579] = 33'd169185942;
        test_addr[1580] = 886;
        test_data[1580] = 33'd3848846976;
        test_addr[1581] = 887;
        test_data[1581] = 33'd2461902253;
        test_addr[1582] = 888;
        test_data[1582] = 33'd2681275051;
        test_addr[1583] = 699;
        test_data[1583] = 33'd7294049884;
        test_addr[1584] = 700;
        test_data[1584] = 33'd1353090612;
        test_addr[1585] = 701;
        test_data[1585] = 33'd3933897631;
        test_addr[1586] = 702;
        test_data[1586] = 33'd5292233811;
        test_addr[1587] = 703;
        test_data[1587] = 33'd5081430845;
        test_addr[1588] = 704;
        test_data[1588] = 33'd5417834559;
        test_addr[1589] = 705;
        test_data[1589] = 33'd1050986732;
        test_addr[1590] = 706;
        test_data[1590] = 33'd6587608098;
        test_addr[1591] = 889;
        test_data[1591] = 33'd6768034894;
        test_addr[1592] = 890;
        test_data[1592] = 33'd1018830267;
        test_addr[1593] = 891;
        test_data[1593] = 33'd4197184161;
        test_addr[1594] = 892;
        test_data[1594] = 33'd1771063249;
        test_addr[1595] = 724;
        test_data[1595] = 33'd3326485598;
        test_addr[1596] = 725;
        test_data[1596] = 33'd6553952119;
        test_addr[1597] = 726;
        test_data[1597] = 33'd4007895896;
        test_addr[1598] = 727;
        test_data[1598] = 33'd2861577116;
        test_addr[1599] = 728;
        test_data[1599] = 33'd2130178182;
        test_addr[1600] = 893;
        test_data[1600] = 33'd2729806528;
        test_addr[1601] = 894;
        test_data[1601] = 33'd1657957379;
        test_addr[1602] = 895;
        test_data[1602] = 33'd1344756801;
        test_addr[1603] = 896;
        test_data[1603] = 33'd1203527177;
        test_addr[1604] = 897;
        test_data[1604] = 33'd1983065030;
        test_addr[1605] = 898;
        test_data[1605] = 33'd4257032184;
        test_addr[1606] = 899;
        test_data[1606] = 33'd2405277136;
        test_addr[1607] = 900;
        test_data[1607] = 33'd3781980178;
        test_addr[1608] = 901;
        test_data[1608] = 33'd6907121802;
        test_addr[1609] = 902;
        test_data[1609] = 33'd8381351077;
        test_addr[1610] = 903;
        test_data[1610] = 33'd4884006566;
        test_addr[1611] = 904;
        test_data[1611] = 33'd2619155067;
        test_addr[1612] = 905;
        test_data[1612] = 33'd5879660817;
        test_addr[1613] = 906;
        test_data[1613] = 33'd1994273950;
        test_addr[1614] = 907;
        test_data[1614] = 33'd1385986733;
        test_addr[1615] = 908;
        test_data[1615] = 33'd214893740;
        test_addr[1616] = 909;
        test_data[1616] = 33'd3200669720;
        test_addr[1617] = 910;
        test_data[1617] = 33'd1125257678;
        test_addr[1618] = 911;
        test_data[1618] = 33'd3639758164;
        test_addr[1619] = 912;
        test_data[1619] = 33'd5821672846;
        test_addr[1620] = 913;
        test_data[1620] = 33'd1701002144;
        test_addr[1621] = 914;
        test_data[1621] = 33'd617611722;
        test_addr[1622] = 915;
        test_data[1622] = 33'd316048180;
        test_addr[1623] = 916;
        test_data[1623] = 33'd8038283157;
        test_addr[1624] = 917;
        test_data[1624] = 33'd347883434;
        test_addr[1625] = 918;
        test_data[1625] = 33'd8395401196;
        test_addr[1626] = 919;
        test_data[1626] = 33'd1993211956;
        test_addr[1627] = 920;
        test_data[1627] = 33'd7592216072;
        test_addr[1628] = 921;
        test_data[1628] = 33'd244390958;
        test_addr[1629] = 922;
        test_data[1629] = 33'd268862713;
        test_addr[1630] = 239;
        test_data[1630] = 33'd3601678559;
        test_addr[1631] = 240;
        test_data[1631] = 33'd272401660;
        test_addr[1632] = 241;
        test_data[1632] = 33'd6487185225;
        test_addr[1633] = 242;
        test_data[1633] = 33'd2915968114;
        test_addr[1634] = 923;
        test_data[1634] = 33'd2554414221;
        test_addr[1635] = 924;
        test_data[1635] = 33'd1164293521;
        test_addr[1636] = 157;
        test_data[1636] = 33'd6917650850;
        test_addr[1637] = 158;
        test_data[1637] = 33'd5997311169;
        test_addr[1638] = 159;
        test_data[1638] = 33'd2928595937;
        test_addr[1639] = 160;
        test_data[1639] = 33'd660917259;
        test_addr[1640] = 161;
        test_data[1640] = 33'd523302279;
        test_addr[1641] = 162;
        test_data[1641] = 33'd6640639342;
        test_addr[1642] = 163;
        test_data[1642] = 33'd6986933559;
        test_addr[1643] = 164;
        test_data[1643] = 33'd8314209422;
        test_addr[1644] = 165;
        test_data[1644] = 33'd117310100;
        test_addr[1645] = 166;
        test_data[1645] = 33'd288407532;
        test_addr[1646] = 167;
        test_data[1646] = 33'd7200750765;
        test_addr[1647] = 168;
        test_data[1647] = 33'd1522146474;
        test_addr[1648] = 169;
        test_data[1648] = 33'd654559525;
        test_addr[1649] = 170;
        test_data[1649] = 33'd574793399;
        test_addr[1650] = 171;
        test_data[1650] = 33'd5465076370;
        test_addr[1651] = 172;
        test_data[1651] = 33'd460255681;
        test_addr[1652] = 173;
        test_data[1652] = 33'd6721134700;
        test_addr[1653] = 174;
        test_data[1653] = 33'd1373713971;
        test_addr[1654] = 175;
        test_data[1654] = 33'd6972805961;
        test_addr[1655] = 176;
        test_data[1655] = 33'd2743796502;
        test_addr[1656] = 177;
        test_data[1656] = 33'd1825087556;
        test_addr[1657] = 178;
        test_data[1657] = 33'd3775849174;
        test_addr[1658] = 925;
        test_data[1658] = 33'd74622926;
        test_addr[1659] = 926;
        test_data[1659] = 33'd2262293352;
        test_addr[1660] = 927;
        test_data[1660] = 33'd5091422264;
        test_addr[1661] = 928;
        test_data[1661] = 33'd3420167902;
        test_addr[1662] = 929;
        test_data[1662] = 33'd940344392;
        test_addr[1663] = 930;
        test_data[1663] = 33'd7763619672;
        test_addr[1664] = 931;
        test_data[1664] = 33'd3103550827;
        test_addr[1665] = 932;
        test_data[1665] = 33'd6968050113;
        test_addr[1666] = 933;
        test_data[1666] = 33'd2511644972;
        test_addr[1667] = 934;
        test_data[1667] = 33'd2823866363;
        test_addr[1668] = 935;
        test_data[1668] = 33'd1717104902;
        test_addr[1669] = 936;
        test_data[1669] = 33'd6079027575;
        test_addr[1670] = 937;
        test_data[1670] = 33'd2203028531;
        test_addr[1671] = 938;
        test_data[1671] = 33'd2400356313;
        test_addr[1672] = 939;
        test_data[1672] = 33'd2075534042;
        test_addr[1673] = 574;
        test_data[1673] = 33'd4557786605;
        test_addr[1674] = 575;
        test_data[1674] = 33'd197152237;
        test_addr[1675] = 940;
        test_data[1675] = 33'd1707455229;
        test_addr[1676] = 941;
        test_data[1676] = 33'd2844599084;
        test_addr[1677] = 942;
        test_data[1677] = 33'd6576089902;
        test_addr[1678] = 943;
        test_data[1678] = 33'd3573192684;
        test_addr[1679] = 944;
        test_data[1679] = 33'd1106836672;
        test_addr[1680] = 945;
        test_data[1680] = 33'd4038263291;
        test_addr[1681] = 946;
        test_data[1681] = 33'd3719653609;
        test_addr[1682] = 947;
        test_data[1682] = 33'd6075128882;
        test_addr[1683] = 948;
        test_data[1683] = 33'd1347233679;
        test_addr[1684] = 949;
        test_data[1684] = 33'd318477808;
        test_addr[1685] = 395;
        test_data[1685] = 33'd2126893221;
        test_addr[1686] = 950;
        test_data[1686] = 33'd1211772756;
        test_addr[1687] = 951;
        test_data[1687] = 33'd4372174755;
        test_addr[1688] = 952;
        test_data[1688] = 33'd3841582932;
        test_addr[1689] = 953;
        test_data[1689] = 33'd1358315614;
        test_addr[1690] = 954;
        test_data[1690] = 33'd3948916793;
        test_addr[1691] = 955;
        test_data[1691] = 33'd976392251;
        test_addr[1692] = 956;
        test_data[1692] = 33'd604891091;
        test_addr[1693] = 957;
        test_data[1693] = 33'd2766494036;
        test_addr[1694] = 649;
        test_data[1694] = 33'd3154846827;
        test_addr[1695] = 650;
        test_data[1695] = 33'd1968337716;
        test_addr[1696] = 651;
        test_data[1696] = 33'd7668884202;
        test_addr[1697] = 652;
        test_data[1697] = 33'd1737322648;
        test_addr[1698] = 653;
        test_data[1698] = 33'd5065262374;
        test_addr[1699] = 654;
        test_data[1699] = 33'd1955032163;
        test_addr[1700] = 655;
        test_data[1700] = 33'd6695552079;
        test_addr[1701] = 656;
        test_data[1701] = 33'd903928419;
        test_addr[1702] = 657;
        test_data[1702] = 33'd4073638024;
        test_addr[1703] = 658;
        test_data[1703] = 33'd420911824;
        test_addr[1704] = 659;
        test_data[1704] = 33'd6318685622;
        test_addr[1705] = 660;
        test_data[1705] = 33'd6345835911;
        test_addr[1706] = 661;
        test_data[1706] = 33'd6344047751;
        test_addr[1707] = 662;
        test_data[1707] = 33'd4771531159;
        test_addr[1708] = 663;
        test_data[1708] = 33'd463783079;
        test_addr[1709] = 664;
        test_data[1709] = 33'd961409848;
        test_addr[1710] = 665;
        test_data[1710] = 33'd5387516243;
        test_addr[1711] = 666;
        test_data[1711] = 33'd3656350260;
        test_addr[1712] = 667;
        test_data[1712] = 33'd7771786512;
        test_addr[1713] = 668;
        test_data[1713] = 33'd2346181448;
        test_addr[1714] = 669;
        test_data[1714] = 33'd3867887075;
        test_addr[1715] = 958;
        test_data[1715] = 33'd6946123739;
        test_addr[1716] = 959;
        test_data[1716] = 33'd1529856229;
        test_addr[1717] = 393;
        test_data[1717] = 33'd2750675278;
        test_addr[1718] = 960;
        test_data[1718] = 33'd1948195766;
        test_addr[1719] = 961;
        test_data[1719] = 33'd2424908381;
        test_addr[1720] = 962;
        test_data[1720] = 33'd1061798646;
        test_addr[1721] = 963;
        test_data[1721] = 33'd116665739;
        test_addr[1722] = 964;
        test_data[1722] = 33'd8317080837;
        test_addr[1723] = 965;
        test_data[1723] = 33'd3248282811;
        test_addr[1724] = 966;
        test_data[1724] = 33'd4155125915;
        test_addr[1725] = 967;
        test_data[1725] = 33'd6733892002;
        test_addr[1726] = 968;
        test_data[1726] = 33'd1749865633;
        test_addr[1727] = 669;
        test_data[1727] = 33'd5238013991;
        test_addr[1728] = 670;
        test_data[1728] = 33'd270318229;
        test_addr[1729] = 671;
        test_data[1729] = 33'd6461600984;
        test_addr[1730] = 969;
        test_data[1730] = 33'd2080802869;
        test_addr[1731] = 970;
        test_data[1731] = 33'd2451347637;
        test_addr[1732] = 971;
        test_data[1732] = 33'd713104100;
        test_addr[1733] = 972;
        test_data[1733] = 33'd3792588729;
        test_addr[1734] = 973;
        test_data[1734] = 33'd1940515451;
        test_addr[1735] = 974;
        test_data[1735] = 33'd947401983;
        test_addr[1736] = 975;
        test_data[1736] = 33'd4850705758;
        test_addr[1737] = 976;
        test_data[1737] = 33'd3450979905;
        test_addr[1738] = 977;
        test_data[1738] = 33'd3853008963;
        test_addr[1739] = 978;
        test_data[1739] = 33'd1522177301;
        test_addr[1740] = 979;
        test_data[1740] = 33'd7432756012;
        test_addr[1741] = 980;
        test_data[1741] = 33'd127768736;
        test_addr[1742] = 981;
        test_data[1742] = 33'd3878255990;
        test_addr[1743] = 982;
        test_data[1743] = 33'd7574700653;
        test_addr[1744] = 983;
        test_data[1744] = 33'd1650122225;
        test_addr[1745] = 984;
        test_data[1745] = 33'd2979938981;
        test_addr[1746] = 985;
        test_data[1746] = 33'd2125246417;
        test_addr[1747] = 986;
        test_data[1747] = 33'd2058768324;
        test_addr[1748] = 987;
        test_data[1748] = 33'd2669326286;
        test_addr[1749] = 988;
        test_data[1749] = 33'd1629806814;
        test_addr[1750] = 989;
        test_data[1750] = 33'd867504778;
        test_addr[1751] = 990;
        test_data[1751] = 33'd4133797271;
        test_addr[1752] = 991;
        test_data[1752] = 33'd4151446151;
        test_addr[1753] = 992;
        test_data[1753] = 33'd112184677;
        test_addr[1754] = 993;
        test_data[1754] = 33'd3829262925;
        test_addr[1755] = 994;
        test_data[1755] = 33'd7265699461;
        test_addr[1756] = 871;
        test_data[1756] = 33'd4813907875;
        test_addr[1757] = 872;
        test_data[1757] = 33'd7805843445;
        test_addr[1758] = 873;
        test_data[1758] = 33'd4514565983;
        test_addr[1759] = 874;
        test_data[1759] = 33'd5895856864;
        test_addr[1760] = 875;
        test_data[1760] = 33'd4043269648;
        test_addr[1761] = 876;
        test_data[1761] = 33'd1362121102;
        test_addr[1762] = 877;
        test_data[1762] = 33'd5886701679;
        test_addr[1763] = 878;
        test_data[1763] = 33'd6064932223;
        test_addr[1764] = 879;
        test_data[1764] = 33'd7030834215;
        test_addr[1765] = 880;
        test_data[1765] = 33'd7776153154;
        test_addr[1766] = 881;
        test_data[1766] = 33'd1205481735;
        test_addr[1767] = 995;
        test_data[1767] = 33'd4310430729;
        test_addr[1768] = 996;
        test_data[1768] = 33'd428556190;
        test_addr[1769] = 997;
        test_data[1769] = 33'd3032800360;
        test_addr[1770] = 998;
        test_data[1770] = 33'd4049855863;
        test_addr[1771] = 999;
        test_data[1771] = 33'd7850279929;
        test_addr[1772] = 1000;
        test_data[1772] = 33'd3487038663;
        test_addr[1773] = 1001;
        test_data[1773] = 33'd3081669374;
        test_addr[1774] = 1002;
        test_data[1774] = 33'd8480044071;
        test_addr[1775] = 1003;
        test_data[1775] = 33'd3486094991;
        test_addr[1776] = 1004;
        test_data[1776] = 33'd3494997726;
        test_addr[1777] = 1005;
        test_data[1777] = 33'd5095303093;
        test_addr[1778] = 1006;
        test_data[1778] = 33'd4197983772;
        test_addr[1779] = 1007;
        test_data[1779] = 33'd492031920;
        test_addr[1780] = 1008;
        test_data[1780] = 33'd2946475741;
        test_addr[1781] = 1009;
        test_data[1781] = 33'd7647611263;
        test_addr[1782] = 1010;
        test_data[1782] = 33'd7135279520;
        test_addr[1783] = 1011;
        test_data[1783] = 33'd5324429110;
        test_addr[1784] = 1012;
        test_data[1784] = 33'd7987172483;
        test_addr[1785] = 1013;
        test_data[1785] = 33'd2547033048;
        test_addr[1786] = 1014;
        test_data[1786] = 33'd1358387716;
        test_addr[1787] = 1015;
        test_data[1787] = 33'd2574971247;
        test_addr[1788] = 1016;
        test_data[1788] = 33'd7822317535;
        test_addr[1789] = 1017;
        test_data[1789] = 33'd4080120458;
        test_addr[1790] = 469;
        test_data[1790] = 33'd8211500379;
        test_addr[1791] = 470;
        test_data[1791] = 33'd3758623902;
        test_addr[1792] = 471;
        test_data[1792] = 33'd4277788026;
        test_addr[1793] = 1018;
        test_data[1793] = 33'd7078932678;
        test_addr[1794] = 1019;
        test_data[1794] = 33'd7102665382;
        test_addr[1795] = 46;
        test_data[1795] = 33'd2921447489;
        test_addr[1796] = 47;
        test_data[1796] = 33'd2684505263;
        test_addr[1797] = 48;
        test_data[1797] = 33'd5077311334;
        test_addr[1798] = 49;
        test_data[1798] = 33'd1390656163;
        test_addr[1799] = 50;
        test_data[1799] = 33'd2480296893;
        test_addr[1800] = 51;
        test_data[1800] = 33'd893530107;
        test_addr[1801] = 52;
        test_data[1801] = 33'd369651485;
        test_addr[1802] = 53;
        test_data[1802] = 33'd2187729913;
        test_addr[1803] = 54;
        test_data[1803] = 33'd5738633716;
        test_addr[1804] = 55;
        test_data[1804] = 33'd7537695275;
        test_addr[1805] = 56;
        test_data[1805] = 33'd5226950425;
        test_addr[1806] = 1020;
        test_data[1806] = 33'd2038773800;
        test_addr[1807] = 1021;
        test_data[1807] = 33'd8421308923;
        test_addr[1808] = 767;
        test_data[1808] = 33'd2928940173;
        test_addr[1809] = 768;
        test_data[1809] = 33'd5836870268;
        test_addr[1810] = 769;
        test_data[1810] = 33'd194866178;
        test_addr[1811] = 770;
        test_data[1811] = 33'd968883625;
        test_addr[1812] = 1022;
        test_data[1812] = 33'd1277705246;
        test_addr[1813] = 1023;
        test_data[1813] = 33'd2086004592;
        test_addr[1814] = 781;
        test_data[1814] = 33'd2253784569;
        test_addr[1815] = 782;
        test_data[1815] = 33'd6400293048;
        test_addr[1816] = 783;
        test_data[1816] = 33'd5896829583;
        test_addr[1817] = 784;
        test_data[1817] = 33'd4324763413;
        test_addr[1818] = 785;
        test_data[1818] = 33'd2691045821;
        test_addr[1819] = 786;
        test_data[1819] = 33'd5513802879;
        test_addr[1820] = 787;
        test_data[1820] = 33'd109264237;
        test_addr[1821] = 788;
        test_data[1821] = 33'd1639691474;
        test_addr[1822] = 789;
        test_data[1822] = 33'd2090407313;
        test_addr[1823] = 790;
        test_data[1823] = 33'd8271951972;
        test_addr[1824] = 791;
        test_data[1824] = 33'd6626636475;
        test_addr[1825] = 792;
        test_data[1825] = 33'd3990341194;
        test_addr[1826] = 793;
        test_data[1826] = 33'd1132372465;
        test_addr[1827] = 794;
        test_data[1827] = 33'd2371798522;
        test_addr[1828] = 795;
        test_data[1828] = 33'd7612960125;
        test_addr[1829] = 796;
        test_data[1829] = 33'd1668815192;
        test_addr[1830] = 797;
        test_data[1830] = 33'd3852826982;
        test_addr[1831] = 798;
        test_data[1831] = 33'd1995026993;
        test_addr[1832] = 799;
        test_data[1832] = 33'd2623245066;
        test_addr[1833] = 800;
        test_data[1833] = 33'd3694851582;
        test_addr[1834] = 801;
        test_data[1834] = 33'd8174766734;
        test_addr[1835] = 802;
        test_data[1835] = 33'd3175044348;
        test_addr[1836] = 803;
        test_data[1836] = 33'd1019510884;
        test_addr[1837] = 804;
        test_data[1837] = 33'd7530848819;
        test_addr[1838] = 805;
        test_data[1838] = 33'd627959300;
        test_addr[1839] = 806;
        test_data[1839] = 33'd3113296974;
        test_addr[1840] = 807;
        test_data[1840] = 33'd1709814211;
        test_addr[1841] = 808;
        test_data[1841] = 33'd3076343433;
        test_addr[1842] = 809;
        test_data[1842] = 33'd4326162914;
        test_addr[1843] = 810;
        test_data[1843] = 33'd5479111943;
        test_addr[1844] = 811;
        test_data[1844] = 33'd7916788073;
        test_addr[1845] = 812;
        test_data[1845] = 33'd2940558418;
        test_addr[1846] = 813;
        test_data[1846] = 33'd1652768965;
        test_addr[1847] = 814;
        test_data[1847] = 33'd1384835374;
        test_addr[1848] = 815;
        test_data[1848] = 33'd8265617095;
        test_addr[1849] = 816;
        test_data[1849] = 33'd96275483;
        test_addr[1850] = 817;
        test_data[1850] = 33'd1666061305;
        test_addr[1851] = 818;
        test_data[1851] = 33'd6803544565;
        test_addr[1852] = 819;
        test_data[1852] = 33'd5962325336;
        test_addr[1853] = 820;
        test_data[1853] = 33'd3676412073;
        test_addr[1854] = 821;
        test_data[1854] = 33'd707615435;
        test_addr[1855] = 822;
        test_data[1855] = 33'd435222120;
        test_addr[1856] = 823;
        test_data[1856] = 33'd7933540958;
        test_addr[1857] = 824;
        test_data[1857] = 33'd1487235996;
        test_addr[1858] = 825;
        test_data[1858] = 33'd276834200;
        test_addr[1859] = 826;
        test_data[1859] = 33'd5883333751;
        test_addr[1860] = 827;
        test_data[1860] = 33'd4776355001;
        test_addr[1861] = 828;
        test_data[1861] = 33'd3353314327;
        test_addr[1862] = 829;
        test_data[1862] = 33'd6277331716;
        test_addr[1863] = 830;
        test_data[1863] = 33'd2929608453;
        test_addr[1864] = 831;
        test_data[1864] = 33'd11545355;
        test_addr[1865] = 832;
        test_data[1865] = 33'd8365330899;
        test_addr[1866] = 833;
        test_data[1866] = 33'd8113452914;
        test_addr[1867] = 834;
        test_data[1867] = 33'd1981444042;
        test_addr[1868] = 835;
        test_data[1868] = 33'd915768184;
        test_addr[1869] = 836;
        test_data[1869] = 33'd2037704408;
        test_addr[1870] = 837;
        test_data[1870] = 33'd6292354088;
        test_addr[1871] = 838;
        test_data[1871] = 33'd924586107;
        test_addr[1872] = 839;
        test_data[1872] = 33'd1862425237;
        test_addr[1873] = 840;
        test_data[1873] = 33'd967968676;
        test_addr[1874] = 841;
        test_data[1874] = 33'd209372675;
        test_addr[1875] = 842;
        test_data[1875] = 33'd4492505524;
        test_addr[1876] = 843;
        test_data[1876] = 33'd4361648510;
        test_addr[1877] = 844;
        test_data[1877] = 33'd4108930760;
        test_addr[1878] = 845;
        test_data[1878] = 33'd3010963361;
        test_addr[1879] = 846;
        test_data[1879] = 33'd1415523632;
        test_addr[1880] = 847;
        test_data[1880] = 33'd2811533726;
        test_addr[1881] = 848;
        test_data[1881] = 33'd6785720582;
        test_addr[1882] = 849;
        test_data[1882] = 33'd5210670346;
        test_addr[1883] = 850;
        test_data[1883] = 33'd3859470178;
        test_addr[1884] = 851;
        test_data[1884] = 33'd8165676555;
        test_addr[1885] = 852;
        test_data[1885] = 33'd3381402385;
        test_addr[1886] = 853;
        test_data[1886] = 33'd2928255153;
        test_addr[1887] = 854;
        test_data[1887] = 33'd4252373770;
        test_addr[1888] = 855;
        test_data[1888] = 33'd3648691299;
        test_addr[1889] = 856;
        test_data[1889] = 33'd3274644583;
        test_addr[1890] = 857;
        test_data[1890] = 33'd2217991288;
        test_addr[1891] = 858;
        test_data[1891] = 33'd6510627754;
        test_addr[1892] = 859;
        test_data[1892] = 33'd7764311278;
        test_addr[1893] = 860;
        test_data[1893] = 33'd2745739626;
        test_addr[1894] = 861;
        test_data[1894] = 33'd1495467381;
        test_addr[1895] = 862;
        test_data[1895] = 33'd3532219985;
        test_addr[1896] = 863;
        test_data[1896] = 33'd2333676472;
        test_addr[1897] = 864;
        test_data[1897] = 33'd7142189735;
        test_addr[1898] = 865;
        test_data[1898] = 33'd6086640944;
        test_addr[1899] = 866;
        test_data[1899] = 33'd284044551;
        test_addr[1900] = 867;
        test_data[1900] = 33'd11628468;
        test_addr[1901] = 868;
        test_data[1901] = 33'd818584801;
        test_addr[1902] = 0;
        test_data[1902] = 33'd812361294;
        test_addr[1903] = 1;
        test_data[1903] = 33'd1897396466;
        test_addr[1904] = 950;
        test_data[1904] = 33'd1211772756;
        test_addr[1905] = 951;
        test_data[1905] = 33'd4481600501;
        test_addr[1906] = 952;
        test_data[1906] = 33'd3841582932;
        test_addr[1907] = 953;
        test_data[1907] = 33'd1358315614;
        test_addr[1908] = 954;
        test_data[1908] = 33'd3948916793;
        test_addr[1909] = 955;
        test_data[1909] = 33'd976392251;
        test_addr[1910] = 956;
        test_data[1910] = 33'd604891091;
        test_addr[1911] = 957;
        test_data[1911] = 33'd2766494036;
        test_addr[1912] = 958;
        test_data[1912] = 33'd2651156443;
        test_addr[1913] = 959;
        test_data[1913] = 33'd6539801529;
        test_addr[1914] = 960;
        test_data[1914] = 33'd6067332930;
        test_addr[1915] = 961;
        test_data[1915] = 33'd5042235847;
        test_addr[1916] = 962;
        test_data[1916] = 33'd1061798646;
        test_addr[1917] = 963;
        test_data[1917] = 33'd6616312562;
        test_addr[1918] = 964;
        test_data[1918] = 33'd6474981332;
        test_addr[1919] = 965;
        test_data[1919] = 33'd3248282811;
        test_addr[1920] = 966;
        test_data[1920] = 33'd4155125915;
        test_addr[1921] = 967;
        test_data[1921] = 33'd6010715935;
        test_addr[1922] = 968;
        test_data[1922] = 33'd1749865633;
        test_addr[1923] = 969;
        test_data[1923] = 33'd4591053368;
        test_addr[1924] = 2;
        test_data[1924] = 33'd1865453439;
        test_addr[1925] = 3;
        test_data[1925] = 33'd1011693257;
        test_addr[1926] = 802;
        test_data[1926] = 33'd4849342358;
        test_addr[1927] = 803;
        test_data[1927] = 33'd7227299843;
        test_addr[1928] = 804;
        test_data[1928] = 33'd3235881523;
        test_addr[1929] = 805;
        test_data[1929] = 33'd627959300;
        test_addr[1930] = 4;
        test_data[1930] = 33'd93557296;
        test_addr[1931] = 5;
        test_data[1931] = 33'd838687445;
        test_addr[1932] = 6;
        test_data[1932] = 33'd5173796523;
        test_addr[1933] = 7;
        test_data[1933] = 33'd3491080214;
        test_addr[1934] = 8;
        test_data[1934] = 33'd1430891515;
        test_addr[1935] = 9;
        test_data[1935] = 33'd1174159001;
        test_addr[1936] = 10;
        test_data[1936] = 33'd1664182063;
        test_addr[1937] = 933;
        test_data[1937] = 33'd2511644972;
        test_addr[1938] = 934;
        test_data[1938] = 33'd2823866363;
        test_addr[1939] = 935;
        test_data[1939] = 33'd5076926062;
        test_addr[1940] = 936;
        test_data[1940] = 33'd7416665667;
        test_addr[1941] = 937;
        test_data[1941] = 33'd8225306977;
        test_addr[1942] = 938;
        test_data[1942] = 33'd4543047013;
        test_addr[1943] = 939;
        test_data[1943] = 33'd2075534042;
        test_addr[1944] = 11;
        test_data[1944] = 33'd773081521;
        test_addr[1945] = 12;
        test_data[1945] = 33'd3296343955;
        test_addr[1946] = 13;
        test_data[1946] = 33'd1476987912;
        test_addr[1947] = 14;
        test_data[1947] = 33'd1747019271;
        test_addr[1948] = 15;
        test_data[1948] = 33'd1389907803;
        test_addr[1949] = 16;
        test_data[1949] = 33'd2995721384;
        test_addr[1950] = 17;
        test_data[1950] = 33'd1707974702;
        test_addr[1951] = 18;
        test_data[1951] = 33'd1571951305;
        test_addr[1952] = 19;
        test_data[1952] = 33'd6095237219;
        test_addr[1953] = 20;
        test_data[1953] = 33'd1223440380;
        test_addr[1954] = 21;
        test_data[1954] = 33'd3366782182;
        test_addr[1955] = 22;
        test_data[1955] = 33'd5698914819;
        test_addr[1956] = 23;
        test_data[1956] = 33'd2361297799;
        test_addr[1957] = 24;
        test_data[1957] = 33'd2711593210;
        test_addr[1958] = 25;
        test_data[1958] = 33'd4002336428;
        test_addr[1959] = 26;
        test_data[1959] = 33'd4291600053;
        test_addr[1960] = 27;
        test_data[1960] = 33'd5269698867;
        test_addr[1961] = 28;
        test_data[1961] = 33'd8248660826;
        test_addr[1962] = 29;
        test_data[1962] = 33'd3331445440;
        test_addr[1963] = 30;
        test_data[1963] = 33'd1741498846;
        test_addr[1964] = 31;
        test_data[1964] = 33'd7375367997;
        test_addr[1965] = 32;
        test_data[1965] = 33'd8046170488;
        test_addr[1966] = 33;
        test_data[1966] = 33'd2359621732;
        test_addr[1967] = 34;
        test_data[1967] = 33'd1887051034;
        test_addr[1968] = 35;
        test_data[1968] = 33'd172683611;
        test_addr[1969] = 36;
        test_data[1969] = 33'd2709550290;
        test_addr[1970] = 37;
        test_data[1970] = 33'd406326701;
        test_addr[1971] = 38;
        test_data[1971] = 33'd300770812;
        test_addr[1972] = 168;
        test_data[1972] = 33'd1522146474;
        test_addr[1973] = 169;
        test_data[1973] = 33'd654559525;
        test_addr[1974] = 170;
        test_data[1974] = 33'd574793399;
        test_addr[1975] = 171;
        test_data[1975] = 33'd1170109074;
        test_addr[1976] = 172;
        test_data[1976] = 33'd4652336758;
        test_addr[1977] = 173;
        test_data[1977] = 33'd2426167404;
        test_addr[1978] = 174;
        test_data[1978] = 33'd1373713971;
        test_addr[1979] = 175;
        test_data[1979] = 33'd7301232615;
        test_addr[1980] = 176;
        test_data[1980] = 33'd2743796502;
        test_addr[1981] = 177;
        test_data[1981] = 33'd1825087556;
        test_addr[1982] = 178;
        test_data[1982] = 33'd3775849174;
        test_addr[1983] = 39;
        test_data[1983] = 33'd1715945728;
        test_addr[1984] = 40;
        test_data[1984] = 33'd4946218338;
        test_addr[1985] = 41;
        test_data[1985] = 33'd2411058451;
        test_addr[1986] = 42;
        test_data[1986] = 33'd2859414406;
        test_addr[1987] = 43;
        test_data[1987] = 33'd389770497;
        test_addr[1988] = 44;
        test_data[1988] = 33'd5205655190;
        test_addr[1989] = 45;
        test_data[1989] = 33'd4991217978;
        test_addr[1990] = 46;
        test_data[1990] = 33'd2921447489;
        test_addr[1991] = 47;
        test_data[1991] = 33'd2684505263;
        test_addr[1992] = 48;
        test_data[1992] = 33'd6403403978;
        test_addr[1993] = 49;
        test_data[1993] = 33'd1390656163;
        test_addr[1994] = 50;
        test_data[1994] = 33'd6594043259;
        test_addr[1995] = 51;
        test_data[1995] = 33'd893530107;
        test_addr[1996] = 52;
        test_data[1996] = 33'd369651485;
        test_addr[1997] = 53;
        test_data[1997] = 33'd2187729913;
        test_addr[1998] = 54;
        test_data[1998] = 33'd1443666420;
        test_addr[1999] = 55;
        test_data[1999] = 33'd4472345505;
        test_addr[2000] = 254;
        test_data[2000] = 33'd6032177246;
        test_addr[2001] = 255;
        test_data[2001] = 33'd5764577843;
        test_addr[2002] = 256;
        test_data[2002] = 33'd2800244347;
        test_addr[2003] = 257;
        test_data[2003] = 33'd3077211561;
        test_addr[2004] = 258;
        test_data[2004] = 33'd5545252506;
        test_addr[2005] = 259;
        test_data[2005] = 33'd791380853;
        test_addr[2006] = 260;
        test_data[2006] = 33'd1766135903;
        test_addr[2007] = 261;
        test_data[2007] = 33'd2250015139;
        test_addr[2008] = 56;
        test_data[2008] = 33'd4390018467;
        test_addr[2009] = 57;
        test_data[2009] = 33'd3485717736;
        test_addr[2010] = 58;
        test_data[2010] = 33'd528146972;
        test_addr[2011] = 59;
        test_data[2011] = 33'd5908691051;
        test_addr[2012] = 60;
        test_data[2012] = 33'd2587167315;
        test_addr[2013] = 61;
        test_data[2013] = 33'd3444518270;
        test_addr[2014] = 1019;
        test_data[2014] = 33'd6183429777;
        test_addr[2015] = 1020;
        test_data[2015] = 33'd2038773800;
        test_addr[2016] = 1021;
        test_data[2016] = 33'd4318012491;
        test_addr[2017] = 1022;
        test_data[2017] = 33'd1277705246;
        test_addr[2018] = 62;
        test_data[2018] = 33'd8084014525;
        test_addr[2019] = 63;
        test_data[2019] = 33'd2080091441;
        test_addr[2020] = 587;
        test_data[2020] = 33'd6178009353;
        test_addr[2021] = 588;
        test_data[2021] = 33'd1568993292;
        test_addr[2022] = 589;
        test_data[2022] = 33'd2295885502;
        test_addr[2023] = 64;
        test_data[2023] = 33'd4280548596;
        test_addr[2024] = 65;
        test_data[2024] = 33'd5537220738;
        test_addr[2025] = 66;
        test_data[2025] = 33'd2358437066;
        test_addr[2026] = 67;
        test_data[2026] = 33'd1974385293;
        test_addr[2027] = 68;
        test_data[2027] = 33'd516941037;
        test_addr[2028] = 69;
        test_data[2028] = 33'd5257542177;
        test_addr[2029] = 70;
        test_data[2029] = 33'd5113604019;
        test_addr[2030] = 30;
        test_data[2030] = 33'd1741498846;
        test_addr[2031] = 71;
        test_data[2031] = 33'd2915912397;
        test_addr[2032] = 72;
        test_data[2032] = 33'd1456092511;
        test_addr[2033] = 73;
        test_data[2033] = 33'd4643893447;
        test_addr[2034] = 74;
        test_data[2034] = 33'd3952396333;
        test_addr[2035] = 75;
        test_data[2035] = 33'd2806077644;
        test_addr[2036] = 76;
        test_data[2036] = 33'd2442953578;
        test_addr[2037] = 77;
        test_data[2037] = 33'd6723729405;
        test_addr[2038] = 78;
        test_data[2038] = 33'd5218852603;
        test_addr[2039] = 79;
        test_data[2039] = 33'd5091210574;
        test_addr[2040] = 80;
        test_data[2040] = 33'd3727744700;
        test_addr[2041] = 81;
        test_data[2041] = 33'd6586299958;
        test_addr[2042] = 82;
        test_data[2042] = 33'd7308771387;
        test_addr[2043] = 83;
        test_data[2043] = 33'd1729932993;
        test_addr[2044] = 84;
        test_data[2044] = 33'd3961820065;
        test_addr[2045] = 320;
        test_data[2045] = 33'd1997760002;
        test_addr[2046] = 321;
        test_data[2046] = 33'd2940510207;
        test_addr[2047] = 322;
        test_data[2047] = 33'd2475824748;
        test_addr[2048] = 323;
        test_data[2048] = 33'd7724311115;
        test_addr[2049] = 324;
        test_data[2049] = 33'd1485894970;
        test_addr[2050] = 325;
        test_data[2050] = 33'd1503820403;
        test_addr[2051] = 326;
        test_data[2051] = 33'd7565750429;
        test_addr[2052] = 327;
        test_data[2052] = 33'd3743832391;
        test_addr[2053] = 328;
        test_data[2053] = 33'd1645146772;
        test_addr[2054] = 329;
        test_data[2054] = 33'd1930974629;
        test_addr[2055] = 330;
        test_data[2055] = 33'd4410547791;
        test_addr[2056] = 331;
        test_data[2056] = 33'd1012710083;
        test_addr[2057] = 332;
        test_data[2057] = 33'd3964024451;
        test_addr[2058] = 85;
        test_data[2058] = 33'd4995722283;
        test_addr[2059] = 86;
        test_data[2059] = 33'd1751965698;
        test_addr[2060] = 87;
        test_data[2060] = 33'd7489491967;
        test_addr[2061] = 88;
        test_data[2061] = 33'd2879312064;
        test_addr[2062] = 89;
        test_data[2062] = 33'd3931536015;
        test_addr[2063] = 90;
        test_data[2063] = 33'd3529518118;
        test_addr[2064] = 91;
        test_data[2064] = 33'd1285586415;
        test_addr[2065] = 92;
        test_data[2065] = 33'd2746581280;
        test_addr[2066] = 24;
        test_data[2066] = 33'd6962127907;
        test_addr[2067] = 25;
        test_data[2067] = 33'd4002336428;
        test_addr[2068] = 26;
        test_data[2068] = 33'd5279877983;
        test_addr[2069] = 27;
        test_data[2069] = 33'd974731571;
        test_addr[2070] = 28;
        test_data[2070] = 33'd3953693530;
        test_addr[2071] = 29;
        test_data[2071] = 33'd3331445440;
        test_addr[2072] = 30;
        test_data[2072] = 33'd7616382774;
        test_addr[2073] = 31;
        test_data[2073] = 33'd6304671681;
        test_addr[2074] = 32;
        test_data[2074] = 33'd3751203192;
        test_addr[2075] = 33;
        test_data[2075] = 33'd2359621732;
        test_addr[2076] = 34;
        test_data[2076] = 33'd1887051034;
        test_addr[2077] = 35;
        test_data[2077] = 33'd172683611;
        test_addr[2078] = 36;
        test_data[2078] = 33'd5241821197;
        test_addr[2079] = 37;
        test_data[2079] = 33'd6899929475;
        test_addr[2080] = 38;
        test_data[2080] = 33'd300770812;
        test_addr[2081] = 39;
        test_data[2081] = 33'd8105083833;
        test_addr[2082] = 40;
        test_data[2082] = 33'd651251042;
        test_addr[2083] = 41;
        test_data[2083] = 33'd7877483466;
        test_addr[2084] = 42;
        test_data[2084] = 33'd6932636219;
        test_addr[2085] = 43;
        test_data[2085] = 33'd389770497;
        test_addr[2086] = 44;
        test_data[2086] = 33'd910687894;
        test_addr[2087] = 45;
        test_data[2087] = 33'd696250682;
        test_addr[2088] = 46;
        test_data[2088] = 33'd2921447489;
        test_addr[2089] = 47;
        test_data[2089] = 33'd2684505263;
        test_addr[2090] = 48;
        test_data[2090] = 33'd2108436682;
        test_addr[2091] = 49;
        test_data[2091] = 33'd1390656163;
        test_addr[2092] = 50;
        test_data[2092] = 33'd2299075963;
        test_addr[2093] = 51;
        test_data[2093] = 33'd893530107;
        test_addr[2094] = 52;
        test_data[2094] = 33'd369651485;
        test_addr[2095] = 53;
        test_data[2095] = 33'd2187729913;
        test_addr[2096] = 54;
        test_data[2096] = 33'd1443666420;
        test_addr[2097] = 55;
        test_data[2097] = 33'd177378209;
        test_addr[2098] = 93;
        test_data[2098] = 33'd3760806334;
        test_addr[2099] = 94;
        test_data[2099] = 33'd8239870588;
        test_addr[2100] = 95;
        test_data[2100] = 33'd4677938537;
        test_addr[2101] = 96;
        test_data[2101] = 33'd5711678601;
        test_addr[2102] = 97;
        test_data[2102] = 33'd8071602235;
        test_addr[2103] = 98;
        test_data[2103] = 33'd5700692492;
        test_addr[2104] = 99;
        test_data[2104] = 33'd5015081651;
        test_addr[2105] = 100;
        test_data[2105] = 33'd1882137235;
        test_addr[2106] = 101;
        test_data[2106] = 33'd2989968304;
        test_addr[2107] = 102;
        test_data[2107] = 33'd3773128195;
        test_addr[2108] = 103;
        test_data[2108] = 33'd1019640399;
        test_addr[2109] = 104;
        test_data[2109] = 33'd4312173855;
        test_addr[2110] = 808;
        test_data[2110] = 33'd3076343433;
        test_addr[2111] = 809;
        test_data[2111] = 33'd31195618;
        test_addr[2112] = 810;
        test_data[2112] = 33'd1184144647;
        test_addr[2113] = 105;
        test_data[2113] = 33'd627517218;
        test_addr[2114] = 956;
        test_data[2114] = 33'd604891091;
        test_addr[2115] = 957;
        test_data[2115] = 33'd6899640757;
        test_addr[2116] = 958;
        test_data[2116] = 33'd2651156443;
        test_addr[2117] = 959;
        test_data[2117] = 33'd2244834233;
        test_addr[2118] = 960;
        test_data[2118] = 33'd1772365634;
        test_addr[2119] = 961;
        test_data[2119] = 33'd747268551;
        test_addr[2120] = 962;
        test_data[2120] = 33'd1061798646;
        test_addr[2121] = 963;
        test_data[2121] = 33'd5981499576;
        test_addr[2122] = 964;
        test_data[2122] = 33'd6370789053;
        test_addr[2123] = 965;
        test_data[2123] = 33'd3248282811;
        test_addr[2124] = 966;
        test_data[2124] = 33'd4155125915;
        test_addr[2125] = 967;
        test_data[2125] = 33'd1715748639;
        test_addr[2126] = 968;
        test_data[2126] = 33'd1749865633;
        test_addr[2127] = 969;
        test_data[2127] = 33'd6961321930;
        test_addr[2128] = 970;
        test_data[2128] = 33'd2451347637;
        test_addr[2129] = 971;
        test_data[2129] = 33'd713104100;
        test_addr[2130] = 972;
        test_data[2130] = 33'd3792588729;
        test_addr[2131] = 973;
        test_data[2131] = 33'd1940515451;
        test_addr[2132] = 974;
        test_data[2132] = 33'd947401983;
        test_addr[2133] = 975;
        test_data[2133] = 33'd8286286889;
        test_addr[2134] = 976;
        test_data[2134] = 33'd3450979905;
        test_addr[2135] = 977;
        test_data[2135] = 33'd3853008963;
        test_addr[2136] = 978;
        test_data[2136] = 33'd1522177301;
        test_addr[2137] = 979;
        test_data[2137] = 33'd3137788716;
        test_addr[2138] = 980;
        test_data[2138] = 33'd127768736;
        test_addr[2139] = 981;
        test_data[2139] = 33'd8156093195;
        test_addr[2140] = 982;
        test_data[2140] = 33'd7579700198;
        test_addr[2141] = 983;
        test_data[2141] = 33'd6895623034;
        test_addr[2142] = 106;
        test_data[2142] = 33'd966105166;
        test_addr[2143] = 107;
        test_data[2143] = 33'd5354004654;
        test_addr[2144] = 108;
        test_data[2144] = 33'd3736950978;
        test_addr[2145] = 109;
        test_data[2145] = 33'd264822472;
        test_addr[2146] = 110;
        test_data[2146] = 33'd7784365863;
        test_addr[2147] = 111;
        test_data[2147] = 33'd645329535;
        test_addr[2148] = 736;
        test_data[2148] = 33'd7838359037;
        test_addr[2149] = 737;
        test_data[2149] = 33'd8580549254;
        test_addr[2150] = 112;
        test_data[2150] = 33'd1815641454;
        test_addr[2151] = 113;
        test_data[2151] = 33'd5775693360;
        test_addr[2152] = 114;
        test_data[2152] = 33'd2554819996;
        test_addr[2153] = 115;
        test_data[2153] = 33'd1121746377;
        test_addr[2154] = 116;
        test_data[2154] = 33'd6144344247;
        test_addr[2155] = 117;
        test_data[2155] = 33'd3966752148;
        test_addr[2156] = 455;
        test_data[2156] = 33'd1395395928;
        test_addr[2157] = 456;
        test_data[2157] = 33'd2711175043;
        test_addr[2158] = 118;
        test_data[2158] = 33'd2078089603;
        test_addr[2159] = 119;
        test_data[2159] = 33'd3539208672;
        test_addr[2160] = 120;
        test_data[2160] = 33'd1032890496;
        test_addr[2161] = 820;
        test_data[2161] = 33'd3676412073;
        test_addr[2162] = 821;
        test_data[2162] = 33'd707615435;
        test_addr[2163] = 822;
        test_data[2163] = 33'd6541126077;
        test_addr[2164] = 823;
        test_data[2164] = 33'd3638573662;
        test_addr[2165] = 824;
        test_data[2165] = 33'd7273569812;
        test_addr[2166] = 825;
        test_data[2166] = 33'd276834200;
        test_addr[2167] = 826;
        test_data[2167] = 33'd1588366455;
        test_addr[2168] = 121;
        test_data[2168] = 33'd557179377;
        test_addr[2169] = 122;
        test_data[2169] = 33'd886188703;
        test_addr[2170] = 123;
        test_data[2170] = 33'd7240569561;
        test_addr[2171] = 124;
        test_data[2171] = 33'd2261534157;
        test_addr[2172] = 125;
        test_data[2172] = 33'd409693294;
        test_addr[2173] = 126;
        test_data[2173] = 33'd717632510;
        test_addr[2174] = 127;
        test_data[2174] = 33'd6166404623;
        test_addr[2175] = 128;
        test_data[2175] = 33'd4085576191;
        test_addr[2176] = 129;
        test_data[2176] = 33'd7898671004;
        test_addr[2177] = 130;
        test_data[2177] = 33'd2760717433;
        test_addr[2178] = 131;
        test_data[2178] = 33'd3219734873;
        test_addr[2179] = 132;
        test_data[2179] = 33'd1457531679;
        test_addr[2180] = 133;
        test_data[2180] = 33'd1165153273;
        test_addr[2181] = 134;
        test_data[2181] = 33'd3496094639;
        test_addr[2182] = 135;
        test_data[2182] = 33'd3470509274;
        test_addr[2183] = 136;
        test_data[2183] = 33'd1366526219;
        test_addr[2184] = 137;
        test_data[2184] = 33'd4277997269;
        test_addr[2185] = 138;
        test_data[2185] = 33'd51940499;
        test_addr[2186] = 341;
        test_data[2186] = 33'd2186863965;
        test_addr[2187] = 139;
        test_data[2187] = 33'd4250352825;
        test_addr[2188] = 140;
        test_data[2188] = 33'd564617519;
        test_addr[2189] = 141;
        test_data[2189] = 33'd485567310;
        test_addr[2190] = 142;
        test_data[2190] = 33'd1458947625;
        test_addr[2191] = 143;
        test_data[2191] = 33'd730436975;
        test_addr[2192] = 144;
        test_data[2192] = 33'd3655464028;
        test_addr[2193] = 145;
        test_data[2193] = 33'd7193443302;
        test_addr[2194] = 146;
        test_data[2194] = 33'd1483917544;
        test_addr[2195] = 147;
        test_data[2195] = 33'd3933851125;
        test_addr[2196] = 148;
        test_data[2196] = 33'd1074274996;
        test_addr[2197] = 149;
        test_data[2197] = 33'd7399210658;
        test_addr[2198] = 150;
        test_data[2198] = 33'd1383869392;
        test_addr[2199] = 151;
        test_data[2199] = 33'd2820628440;
        test_addr[2200] = 152;
        test_data[2200] = 33'd1326911526;
        test_addr[2201] = 153;
        test_data[2201] = 33'd327985978;
        test_addr[2202] = 39;
        test_data[2202] = 33'd6189278946;
        test_addr[2203] = 40;
        test_data[2203] = 33'd651251042;
        test_addr[2204] = 154;
        test_data[2204] = 33'd412214464;
        test_addr[2205] = 155;
        test_data[2205] = 33'd3182442945;
        test_addr[2206] = 156;
        test_data[2206] = 33'd6026486349;
        test_addr[2207] = 157;
        test_data[2207] = 33'd7228207125;
        test_addr[2208] = 158;
        test_data[2208] = 33'd1702343873;
        test_addr[2209] = 159;
        test_data[2209] = 33'd5134030771;
        test_addr[2210] = 160;
        test_data[2210] = 33'd660917259;
        test_addr[2211] = 161;
        test_data[2211] = 33'd523302279;
        test_addr[2212] = 162;
        test_data[2212] = 33'd5482055859;
        test_addr[2213] = 163;
        test_data[2213] = 33'd4864053908;
        test_addr[2214] = 164;
        test_data[2214] = 33'd4019242126;
        test_addr[2215] = 165;
        test_data[2215] = 33'd117310100;
        test_addr[2216] = 166;
        test_data[2216] = 33'd288407532;
        test_addr[2217] = 167;
        test_data[2217] = 33'd2905783469;
        test_addr[2218] = 168;
        test_data[2218] = 33'd5268165974;
        test_addr[2219] = 169;
        test_data[2219] = 33'd654559525;
        test_addr[2220] = 170;
        test_data[2220] = 33'd574793399;
        test_addr[2221] = 416;
        test_data[2221] = 33'd1219202730;
        test_addr[2222] = 417;
        test_data[2222] = 33'd6306349889;
        test_addr[2223] = 418;
        test_data[2223] = 33'd8096293744;
        test_addr[2224] = 419;
        test_data[2224] = 33'd7494297738;
        test_addr[2225] = 420;
        test_data[2225] = 33'd3910550806;
        test_addr[2226] = 171;
        test_data[2226] = 33'd1170109074;
        test_addr[2227] = 172;
        test_data[2227] = 33'd357369462;
        test_addr[2228] = 173;
        test_data[2228] = 33'd2426167404;
        test_addr[2229] = 174;
        test_data[2229] = 33'd1373713971;
        test_addr[2230] = 175;
        test_data[2230] = 33'd3006265319;
        test_addr[2231] = 176;
        test_data[2231] = 33'd2743796502;
        test_addr[2232] = 177;
        test_data[2232] = 33'd7698299525;
        test_addr[2233] = 178;
        test_data[2233] = 33'd3775849174;
        test_addr[2234] = 179;
        test_data[2234] = 33'd1928357839;
        test_addr[2235] = 180;
        test_data[2235] = 33'd5074585252;
        test_addr[2236] = 181;
        test_data[2236] = 33'd1495804814;
        test_addr[2237] = 182;
        test_data[2237] = 33'd557477877;
        test_addr[2238] = 183;
        test_data[2238] = 33'd4790449638;
        test_addr[2239] = 184;
        test_data[2239] = 33'd3207147966;
        test_addr[2240] = 185;
        test_data[2240] = 33'd76388760;
        test_addr[2241] = 186;
        test_data[2241] = 33'd3665623001;
        test_addr[2242] = 187;
        test_data[2242] = 33'd800185981;
        test_addr[2243] = 484;
        test_data[2243] = 33'd4269737784;
        test_addr[2244] = 485;
        test_data[2244] = 33'd3345226134;
        test_addr[2245] = 486;
        test_data[2245] = 33'd1324217527;
        test_addr[2246] = 487;
        test_data[2246] = 33'd459174225;
        test_addr[2247] = 488;
        test_data[2247] = 33'd471720366;
        test_addr[2248] = 489;
        test_data[2248] = 33'd1491360199;
        test_addr[2249] = 490;
        test_data[2249] = 33'd3214783106;
        test_addr[2250] = 491;
        test_data[2250] = 33'd7796594285;
        test_addr[2251] = 492;
        test_data[2251] = 33'd7671396072;
        test_addr[2252] = 493;
        test_data[2252] = 33'd5174705254;
        test_addr[2253] = 494;
        test_data[2253] = 33'd821347042;
        test_addr[2254] = 495;
        test_data[2254] = 33'd2117462048;
        test_addr[2255] = 496;
        test_data[2255] = 33'd3581785694;
        test_addr[2256] = 497;
        test_data[2256] = 33'd1177368502;
        test_addr[2257] = 498;
        test_data[2257] = 33'd3822144455;
        test_addr[2258] = 499;
        test_data[2258] = 33'd8292067615;
        test_addr[2259] = 500;
        test_data[2259] = 33'd8017666951;
        test_addr[2260] = 501;
        test_data[2260] = 33'd595715914;
        test_addr[2261] = 502;
        test_data[2261] = 33'd1457378795;
        test_addr[2262] = 503;
        test_data[2262] = 33'd4308773176;
        test_addr[2263] = 504;
        test_data[2263] = 33'd2586581290;
        test_addr[2264] = 505;
        test_data[2264] = 33'd2328699311;
        test_addr[2265] = 188;
        test_data[2265] = 33'd3517196253;
        test_addr[2266] = 189;
        test_data[2266] = 33'd5571962890;
        test_addr[2267] = 190;
        test_data[2267] = 33'd5367196838;
        test_addr[2268] = 191;
        test_data[2268] = 33'd2734067735;
        test_addr[2269] = 192;
        test_data[2269] = 33'd1416109369;
        test_addr[2270] = 193;
        test_data[2270] = 33'd2663489104;
        test_addr[2271] = 194;
        test_data[2271] = 33'd7313564897;
        test_addr[2272] = 195;
        test_data[2272] = 33'd284779812;
        test_addr[2273] = 196;
        test_data[2273] = 33'd4510715005;
        test_addr[2274] = 481;
        test_data[2274] = 33'd3956236381;
        test_addr[2275] = 482;
        test_data[2275] = 33'd3069633443;
        test_addr[2276] = 483;
        test_data[2276] = 33'd2649187208;
        test_addr[2277] = 484;
        test_data[2277] = 33'd4269737784;
        test_addr[2278] = 485;
        test_data[2278] = 33'd3345226134;
        test_addr[2279] = 486;
        test_data[2279] = 33'd1324217527;
        test_addr[2280] = 487;
        test_data[2280] = 33'd459174225;
        test_addr[2281] = 488;
        test_data[2281] = 33'd4317680627;
        test_addr[2282] = 489;
        test_data[2282] = 33'd8245788042;
        test_addr[2283] = 490;
        test_data[2283] = 33'd3214783106;
        test_addr[2284] = 491;
        test_data[2284] = 33'd3501626989;
        test_addr[2285] = 492;
        test_data[2285] = 33'd6104632453;
        test_addr[2286] = 493;
        test_data[2286] = 33'd879737958;
        test_addr[2287] = 494;
        test_data[2287] = 33'd821347042;
        test_addr[2288] = 495;
        test_data[2288] = 33'd2117462048;
        test_addr[2289] = 496;
        test_data[2289] = 33'd3581785694;
        test_addr[2290] = 497;
        test_data[2290] = 33'd1177368502;
        test_addr[2291] = 498;
        test_data[2291] = 33'd3822144455;
        test_addr[2292] = 197;
        test_data[2292] = 33'd2750204444;
        test_addr[2293] = 198;
        test_data[2293] = 33'd4368154383;
        test_addr[2294] = 352;
        test_data[2294] = 33'd3547444809;
        test_addr[2295] = 353;
        test_data[2295] = 33'd3374898901;
        test_addr[2296] = 354;
        test_data[2296] = 33'd701425537;
        test_addr[2297] = 355;
        test_data[2297] = 33'd5759146962;
        test_addr[2298] = 356;
        test_data[2298] = 33'd2020066253;
        test_addr[2299] = 357;
        test_data[2299] = 33'd6984410994;
        test_addr[2300] = 358;
        test_data[2300] = 33'd2161533557;
        test_addr[2301] = 359;
        test_data[2301] = 33'd2495672481;
        test_addr[2302] = 360;
        test_data[2302] = 33'd1452465810;
        test_addr[2303] = 361;
        test_data[2303] = 33'd8291375727;
        test_addr[2304] = 362;
        test_data[2304] = 33'd2841382309;
        test_addr[2305] = 363;
        test_data[2305] = 33'd7155771971;
        test_addr[2306] = 364;
        test_data[2306] = 33'd6100967515;
        test_addr[2307] = 365;
        test_data[2307] = 33'd7622933226;
        test_addr[2308] = 366;
        test_data[2308] = 33'd3707227066;
        test_addr[2309] = 367;
        test_data[2309] = 33'd1471019555;
        test_addr[2310] = 368;
        test_data[2310] = 33'd6199346088;
        test_addr[2311] = 199;
        test_data[2311] = 33'd2378011170;
        test_addr[2312] = 200;
        test_data[2312] = 33'd4250933843;
        test_addr[2313] = 201;
        test_data[2313] = 33'd3717101577;
        test_addr[2314] = 202;
        test_data[2314] = 33'd7187890079;
        test_addr[2315] = 203;
        test_data[2315] = 33'd998547257;
        test_addr[2316] = 578;
        test_data[2316] = 33'd741309116;
        test_addr[2317] = 579;
        test_data[2317] = 33'd3286825499;
        test_addr[2318] = 580;
        test_data[2318] = 33'd4671529079;
        test_addr[2319] = 204;
        test_data[2319] = 33'd2620591812;
        test_addr[2320] = 231;
        test_data[2320] = 33'd6574837166;
        test_addr[2321] = 232;
        test_data[2321] = 33'd1883974499;
        test_addr[2322] = 233;
        test_data[2322] = 33'd2957499205;
        test_addr[2323] = 234;
        test_data[2323] = 33'd4644950679;
        test_addr[2324] = 235;
        test_data[2324] = 33'd3439453128;
        test_addr[2325] = 236;
        test_data[2325] = 33'd4371450794;
        test_addr[2326] = 237;
        test_data[2326] = 33'd1383156410;
        test_addr[2327] = 238;
        test_data[2327] = 33'd736219013;
        test_addr[2328] = 239;
        test_data[2328] = 33'd8467273735;
        test_addr[2329] = 240;
        test_data[2329] = 33'd6109278689;
        test_addr[2330] = 241;
        test_data[2330] = 33'd5564965614;
        test_addr[2331] = 205;
        test_data[2331] = 33'd2964469971;
        test_addr[2332] = 206;
        test_data[2332] = 33'd1330142089;
        test_addr[2333] = 207;
        test_data[2333] = 33'd155196010;
        test_addr[2334] = 208;
        test_data[2334] = 33'd2056872922;
        test_addr[2335] = 209;
        test_data[2335] = 33'd8491703780;
        test_addr[2336] = 210;
        test_data[2336] = 33'd3137301976;
        test_addr[2337] = 211;
        test_data[2337] = 33'd2875926310;
        test_addr[2338] = 212;
        test_data[2338] = 33'd5687235698;
        test_addr[2339] = 213;
        test_data[2339] = 33'd2959424098;
        test_addr[2340] = 214;
        test_data[2340] = 33'd8062353645;
        test_addr[2341] = 215;
        test_data[2341] = 33'd6282179165;
        test_addr[2342] = 216;
        test_data[2342] = 33'd4396846135;
        test_addr[2343] = 217;
        test_data[2343] = 33'd1119239002;
        test_addr[2344] = 218;
        test_data[2344] = 33'd6690619681;
        test_addr[2345] = 219;
        test_data[2345] = 33'd6886327984;
        test_addr[2346] = 220;
        test_data[2346] = 33'd5954410058;
        test_addr[2347] = 221;
        test_data[2347] = 33'd1801818893;
        test_addr[2348] = 222;
        test_data[2348] = 33'd727510908;
        test_addr[2349] = 223;
        test_data[2349] = 33'd4769279352;
        test_addr[2350] = 224;
        test_data[2350] = 33'd5690711169;
        test_addr[2351] = 225;
        test_data[2351] = 33'd3019194714;
        test_addr[2352] = 226;
        test_data[2352] = 33'd4281849382;
        test_addr[2353] = 227;
        test_data[2353] = 33'd1667423717;
        test_addr[2354] = 228;
        test_data[2354] = 33'd46709375;
        test_addr[2355] = 229;
        test_data[2355] = 33'd5942086265;
        test_addr[2356] = 230;
        test_data[2356] = 33'd3332009274;
        test_addr[2357] = 231;
        test_data[2357] = 33'd5939931659;
        test_addr[2358] = 232;
        test_data[2358] = 33'd1883974499;
        test_addr[2359] = 233;
        test_data[2359] = 33'd2957499205;
        test_addr[2360] = 234;
        test_data[2360] = 33'd349983383;
        test_addr[2361] = 235;
        test_data[2361] = 33'd3439453128;
        test_addr[2362] = 236;
        test_data[2362] = 33'd76483498;
        test_addr[2363] = 237;
        test_data[2363] = 33'd6291453718;
        test_addr[2364] = 238;
        test_data[2364] = 33'd736219013;
        test_addr[2365] = 239;
        test_data[2365] = 33'd5347317684;
        test_addr[2366] = 240;
        test_data[2366] = 33'd1814311393;
        test_addr[2367] = 241;
        test_data[2367] = 33'd4546627463;
        test_addr[2368] = 391;
        test_data[2368] = 33'd2712963902;
        test_addr[2369] = 392;
        test_data[2369] = 33'd1088256129;
        test_addr[2370] = 393;
        test_data[2370] = 33'd2750675278;
        test_addr[2371] = 394;
        test_data[2371] = 33'd862789604;
        test_addr[2372] = 395;
        test_data[2372] = 33'd2126893221;
        test_addr[2373] = 396;
        test_data[2373] = 33'd4286897536;
        test_addr[2374] = 397;
        test_data[2374] = 33'd1575257700;
        test_addr[2375] = 398;
        test_data[2375] = 33'd3564413496;
        test_addr[2376] = 399;
        test_data[2376] = 33'd4053828411;
        test_addr[2377] = 400;
        test_data[2377] = 33'd523664291;
        test_addr[2378] = 401;
        test_data[2378] = 33'd1851728206;
        test_addr[2379] = 402;
        test_data[2379] = 33'd3042682872;
        test_addr[2380] = 403;
        test_data[2380] = 33'd8385715967;
        test_addr[2381] = 404;
        test_data[2381] = 33'd478746838;
        test_addr[2382] = 405;
        test_data[2382] = 33'd1215199985;
        test_addr[2383] = 406;
        test_data[2383] = 33'd6371290897;
        test_addr[2384] = 242;
        test_data[2384] = 33'd2915968114;
        test_addr[2385] = 243;
        test_data[2385] = 33'd2004278974;
        test_addr[2386] = 244;
        test_data[2386] = 33'd1146573824;
        test_addr[2387] = 177;
        test_data[2387] = 33'd3403332229;
        test_addr[2388] = 178;
        test_data[2388] = 33'd3775849174;
        test_addr[2389] = 179;
        test_data[2389] = 33'd1928357839;
        test_addr[2390] = 180;
        test_data[2390] = 33'd779617956;
        test_addr[2391] = 181;
        test_data[2391] = 33'd1495804814;
        test_addr[2392] = 182;
        test_data[2392] = 33'd557477877;
        test_addr[2393] = 183;
        test_data[2393] = 33'd495482342;
        test_addr[2394] = 184;
        test_data[2394] = 33'd3207147966;
        test_addr[2395] = 185;
        test_data[2395] = 33'd7899109505;
        test_addr[2396] = 186;
        test_data[2396] = 33'd3665623001;
        test_addr[2397] = 187;
        test_data[2397] = 33'd5112573254;
        test_addr[2398] = 188;
        test_data[2398] = 33'd7243830831;
        test_addr[2399] = 189;
        test_data[2399] = 33'd4791195586;
        test_addr[2400] = 190;
        test_data[2400] = 33'd4652936057;
        test_addr[2401] = 191;
        test_data[2401] = 33'd2734067735;
        test_addr[2402] = 192;
        test_data[2402] = 33'd6725015467;
        test_addr[2403] = 193;
        test_data[2403] = 33'd2663489104;
        test_addr[2404] = 194;
        test_data[2404] = 33'd6387814685;
        test_addr[2405] = 195;
        test_data[2405] = 33'd284779812;
        test_addr[2406] = 196;
        test_data[2406] = 33'd215747709;
        test_addr[2407] = 197;
        test_data[2407] = 33'd2750204444;
        test_addr[2408] = 198;
        test_data[2408] = 33'd73187087;
        test_addr[2409] = 199;
        test_data[2409] = 33'd2378011170;
        test_addr[2410] = 200;
        test_data[2410] = 33'd4250933843;
        test_addr[2411] = 201;
        test_data[2411] = 33'd3717101577;
        test_addr[2412] = 202;
        test_data[2412] = 33'd5296697618;
        test_addr[2413] = 203;
        test_data[2413] = 33'd7457756013;
        test_addr[2414] = 204;
        test_data[2414] = 33'd2620591812;
        test_addr[2415] = 205;
        test_data[2415] = 33'd8106998235;
        test_addr[2416] = 206;
        test_data[2416] = 33'd1330142089;
        test_addr[2417] = 207;
        test_data[2417] = 33'd155196010;
        test_addr[2418] = 208;
        test_data[2418] = 33'd2056872922;
        test_addr[2419] = 209;
        test_data[2419] = 33'd4196736484;
        test_addr[2420] = 210;
        test_data[2420] = 33'd3137301976;
        test_addr[2421] = 211;
        test_data[2421] = 33'd2875926310;
        test_addr[2422] = 212;
        test_data[2422] = 33'd1392268402;
        test_addr[2423] = 213;
        test_data[2423] = 33'd2959424098;
        test_addr[2424] = 214;
        test_data[2424] = 33'd3767386349;
        test_addr[2425] = 215;
        test_data[2425] = 33'd5228041519;
        test_addr[2426] = 216;
        test_data[2426] = 33'd101878839;
        test_addr[2427] = 217;
        test_data[2427] = 33'd4873599768;
        test_addr[2428] = 218;
        test_data[2428] = 33'd6992534742;
        test_addr[2429] = 219;
        test_data[2429] = 33'd2591360688;
        test_addr[2430] = 220;
        test_data[2430] = 33'd4719737456;
        test_addr[2431] = 221;
        test_data[2431] = 33'd4997519548;
        test_addr[2432] = 245;
        test_data[2432] = 33'd6821333162;
        test_addr[2433] = 246;
        test_data[2433] = 33'd348319993;
        test_addr[2434] = 247;
        test_data[2434] = 33'd1238703566;
        test_addr[2435] = 248;
        test_data[2435] = 33'd5520457115;
        test_addr[2436] = 249;
        test_data[2436] = 33'd8192841855;
        test_addr[2437] = 250;
        test_data[2437] = 33'd8431532221;
        test_addr[2438] = 251;
        test_data[2438] = 33'd4785832810;
        test_addr[2439] = 252;
        test_data[2439] = 33'd3216848485;
        test_addr[2440] = 253;
        test_data[2440] = 33'd6417022567;
        test_addr[2441] = 254;
        test_data[2441] = 33'd8120685563;
        test_addr[2442] = 255;
        test_data[2442] = 33'd1469610547;
        test_addr[2443] = 106;
        test_data[2443] = 33'd5074592373;
        test_addr[2444] = 107;
        test_data[2444] = 33'd1059037358;
        test_addr[2445] = 108;
        test_data[2445] = 33'd3736950978;
        test_addr[2446] = 109;
        test_data[2446] = 33'd264822472;
        test_addr[2447] = 110;
        test_data[2447] = 33'd3489398567;
        test_addr[2448] = 111;
        test_data[2448] = 33'd7103898731;
        test_addr[2449] = 112;
        test_data[2449] = 33'd1815641454;
        test_addr[2450] = 113;
        test_data[2450] = 33'd4316750137;
        test_addr[2451] = 114;
        test_data[2451] = 33'd2554819996;
        test_addr[2452] = 115;
        test_data[2452] = 33'd1121746377;
        test_addr[2453] = 116;
        test_data[2453] = 33'd1849376951;
        test_addr[2454] = 117;
        test_data[2454] = 33'd3966752148;
        test_addr[2455] = 118;
        test_data[2455] = 33'd4927413122;
        test_addr[2456] = 256;
        test_data[2456] = 33'd2800244347;
        test_addr[2457] = 257;
        test_data[2457] = 33'd7220461089;
        test_addr[2458] = 258;
        test_data[2458] = 33'd7800975412;
        test_addr[2459] = 259;
        test_data[2459] = 33'd8093541333;
        test_addr[2460] = 260;
        test_data[2460] = 33'd1766135903;
        test_addr[2461] = 261;
        test_data[2461] = 33'd7835078233;
        test_addr[2462] = 262;
        test_data[2462] = 33'd3746748856;
        test_addr[2463] = 263;
        test_data[2463] = 33'd2114950029;
        test_addr[2464] = 264;
        test_data[2464] = 33'd1735708751;
        test_addr[2465] = 265;
        test_data[2465] = 33'd5411453991;
        test_addr[2466] = 266;
        test_data[2466] = 33'd8470576713;
        test_addr[2467] = 267;
        test_data[2467] = 33'd2041453479;
        test_addr[2468] = 268;
        test_data[2468] = 33'd7342953263;
        test_addr[2469] = 269;
        test_data[2469] = 33'd3034594309;
        test_addr[2470] = 847;
        test_data[2470] = 33'd5756011311;
        test_addr[2471] = 848;
        test_data[2471] = 33'd2490753286;
        test_addr[2472] = 849;
        test_data[2472] = 33'd915703050;
        test_addr[2473] = 850;
        test_data[2473] = 33'd3859470178;
        test_addr[2474] = 851;
        test_data[2474] = 33'd3870709259;
        test_addr[2475] = 852;
        test_data[2475] = 33'd3381402385;
        test_addr[2476] = 270;
        test_data[2476] = 33'd3506364173;
        test_addr[2477] = 271;
        test_data[2477] = 33'd2102264294;
        test_addr[2478] = 272;
        test_data[2478] = 33'd5343571337;
        test_addr[2479] = 273;
        test_data[2479] = 33'd2319337381;
        test_addr[2480] = 274;
        test_data[2480] = 33'd1669442267;
        test_addr[2481] = 275;
        test_data[2481] = 33'd3413279259;
        test_addr[2482] = 276;
        test_data[2482] = 33'd5996466521;
        test_addr[2483] = 277;
        test_data[2483] = 33'd2701917713;
        test_addr[2484] = 278;
        test_data[2484] = 33'd2430218657;
        test_addr[2485] = 279;
        test_data[2485] = 33'd1180435179;
        test_addr[2486] = 280;
        test_data[2486] = 33'd2884868618;
        test_addr[2487] = 281;
        test_data[2487] = 33'd569891205;
        test_addr[2488] = 282;
        test_data[2488] = 33'd5945865297;
        test_addr[2489] = 283;
        test_data[2489] = 33'd117234014;
        test_addr[2490] = 284;
        test_data[2490] = 33'd3405728430;
        test_addr[2491] = 285;
        test_data[2491] = 33'd7964635605;
        test_addr[2492] = 286;
        test_data[2492] = 33'd775168527;
        test_addr[2493] = 287;
        test_data[2493] = 33'd6282931027;
        test_addr[2494] = 288;
        test_data[2494] = 33'd1151781196;
        test_addr[2495] = 886;
        test_data[2495] = 33'd7203846115;
        test_addr[2496] = 289;
        test_data[2496] = 33'd6081312203;
        test_addr[2497] = 164;
        test_data[2497] = 33'd4019242126;
        test_addr[2498] = 165;
        test_data[2498] = 33'd6389647514;
        test_addr[2499] = 166;
        test_data[2499] = 33'd7599949664;
        test_addr[2500] = 167;
        test_data[2500] = 33'd7824053807;
        test_addr[2501] = 168;
        test_data[2501] = 33'd973198678;
        test_addr[2502] = 169;
        test_data[2502] = 33'd8305977980;
        test_addr[2503] = 170;
        test_data[2503] = 33'd5630515611;
        test_addr[2504] = 171;
        test_data[2504] = 33'd1170109074;
        test_addr[2505] = 172;
        test_data[2505] = 33'd7838710061;
        test_addr[2506] = 173;
        test_data[2506] = 33'd2426167404;
        test_addr[2507] = 174;
        test_data[2507] = 33'd1373713971;
        test_addr[2508] = 175;
        test_data[2508] = 33'd3006265319;
        test_addr[2509] = 290;
        test_data[2509] = 33'd967556824;
        test_addr[2510] = 291;
        test_data[2510] = 33'd7870853172;
        test_addr[2511] = 292;
        test_data[2511] = 33'd1426556317;
        test_addr[2512] = 293;
        test_data[2512] = 33'd688835068;
        test_addr[2513] = 294;
        test_data[2513] = 33'd5913274493;
        test_addr[2514] = 295;
        test_data[2514] = 33'd2347942712;
        test_addr[2515] = 296;
        test_data[2515] = 33'd1233127960;
        test_addr[2516] = 297;
        test_data[2516] = 33'd3955483560;
        test_addr[2517] = 298;
        test_data[2517] = 33'd7226975756;
        test_addr[2518] = 299;
        test_data[2518] = 33'd5886409493;
        test_addr[2519] = 300;
        test_data[2519] = 33'd1320963640;
        test_addr[2520] = 301;
        test_data[2520] = 33'd2660948838;
        test_addr[2521] = 302;
        test_data[2521] = 33'd7013297358;
        test_addr[2522] = 303;
        test_data[2522] = 33'd5960544866;
        test_addr[2523] = 304;
        test_data[2523] = 33'd7841227820;
        test_addr[2524] = 305;
        test_data[2524] = 33'd4704313432;
        test_addr[2525] = 306;
        test_data[2525] = 33'd621355406;
        test_addr[2526] = 307;
        test_data[2526] = 33'd299096324;
        test_addr[2527] = 308;
        test_data[2527] = 33'd3983220710;
        test_addr[2528] = 309;
        test_data[2528] = 33'd7647197850;
        test_addr[2529] = 310;
        test_data[2529] = 33'd4071754507;
        test_addr[2530] = 311;
        test_data[2530] = 33'd3158301700;
        test_addr[2531] = 312;
        test_data[2531] = 33'd3915746261;
        test_addr[2532] = 313;
        test_data[2532] = 33'd494624070;
        test_addr[2533] = 314;
        test_data[2533] = 33'd8576854580;
        test_addr[2534] = 776;
        test_data[2534] = 33'd2515051088;
        test_addr[2535] = 777;
        test_data[2535] = 33'd5166333867;
        test_addr[2536] = 778;
        test_data[2536] = 33'd4928696111;
        test_addr[2537] = 779;
        test_data[2537] = 33'd5025128489;
        test_addr[2538] = 780;
        test_data[2538] = 33'd7602194058;
        test_addr[2539] = 781;
        test_data[2539] = 33'd2253784569;
        test_addr[2540] = 782;
        test_data[2540] = 33'd2105325752;
        test_addr[2541] = 783;
        test_data[2541] = 33'd6846852221;
        test_addr[2542] = 784;
        test_data[2542] = 33'd29796117;
        test_addr[2543] = 315;
        test_data[2543] = 33'd1132837972;
        test_addr[2544] = 316;
        test_data[2544] = 33'd2860683439;
        test_addr[2545] = 317;
        test_data[2545] = 33'd566819812;
        test_addr[2546] = 318;
        test_data[2546] = 33'd3655450011;
        test_addr[2547] = 319;
        test_data[2547] = 33'd8536808778;
        test_addr[2548] = 320;
        test_data[2548] = 33'd6195849814;
        test_addr[2549] = 321;
        test_data[2549] = 33'd5865774354;
        test_addr[2550] = 322;
        test_data[2550] = 33'd2475824748;
        test_addr[2551] = 323;
        test_data[2551] = 33'd3429343819;
        test_addr[2552] = 324;
        test_data[2552] = 33'd1485894970;
        test_addr[2553] = 325;
        test_data[2553] = 33'd6257551620;
        test_addr[2554] = 326;
        test_data[2554] = 33'd6052692756;
        test_addr[2555] = 327;
        test_data[2555] = 33'd3743832391;
        test_addr[2556] = 328;
        test_data[2556] = 33'd1645146772;
        test_addr[2557] = 329;
        test_data[2557] = 33'd8569911227;
        test_addr[2558] = 330;
        test_data[2558] = 33'd5496849686;
        test_addr[2559] = 331;
        test_data[2559] = 33'd4733107250;
        test_addr[2560] = 332;
        test_data[2560] = 33'd6262637485;
        test_addr[2561] = 333;
        test_data[2561] = 33'd1019459317;
        test_addr[2562] = 334;
        test_data[2562] = 33'd1631873129;
        test_addr[2563] = 335;
        test_data[2563] = 33'd5879008937;
        test_addr[2564] = 336;
        test_data[2564] = 33'd6963134911;
        test_addr[2565] = 337;
        test_data[2565] = 33'd190701906;
        test_addr[2566] = 338;
        test_data[2566] = 33'd2063414812;
        test_addr[2567] = 339;
        test_data[2567] = 33'd2384267827;
        test_addr[2568] = 340;
        test_data[2568] = 33'd4413043891;
        test_addr[2569] = 341;
        test_data[2569] = 33'd2186863965;
        test_addr[2570] = 342;
        test_data[2570] = 33'd4078357046;
        test_addr[2571] = 343;
        test_data[2571] = 33'd3214848827;
        test_addr[2572] = 344;
        test_data[2572] = 33'd3796226835;
        test_addr[2573] = 345;
        test_data[2573] = 33'd1689992503;
        test_addr[2574] = 346;
        test_data[2574] = 33'd3177845839;
        test_addr[2575] = 347;
        test_data[2575] = 33'd1349350927;
        test_addr[2576] = 837;
        test_data[2576] = 33'd1997386792;
        test_addr[2577] = 838;
        test_data[2577] = 33'd924586107;
        test_addr[2578] = 839;
        test_data[2578] = 33'd1862425237;
        test_addr[2579] = 840;
        test_data[2579] = 33'd967968676;
        test_addr[2580] = 841;
        test_data[2580] = 33'd209372675;
        test_addr[2581] = 842;
        test_data[2581] = 33'd197538228;
        test_addr[2582] = 843;
        test_data[2582] = 33'd66681214;
        test_addr[2583] = 844;
        test_data[2583] = 33'd4108930760;
        test_addr[2584] = 845;
        test_data[2584] = 33'd3010963361;
        test_addr[2585] = 846;
        test_data[2585] = 33'd1415523632;
        test_addr[2586] = 348;
        test_data[2586] = 33'd1905133107;
        test_addr[2587] = 315;
        test_data[2587] = 33'd6222138684;
        test_addr[2588] = 316;
        test_data[2588] = 33'd2860683439;
        test_addr[2589] = 317;
        test_data[2589] = 33'd566819812;
        test_addr[2590] = 318;
        test_data[2590] = 33'd3655450011;
        test_addr[2591] = 319;
        test_data[2591] = 33'd6044180141;
        test_addr[2592] = 320;
        test_data[2592] = 33'd1900882518;
        test_addr[2593] = 321;
        test_data[2593] = 33'd1570807058;
        test_addr[2594] = 349;
        test_data[2594] = 33'd3684863624;
        test_addr[2595] = 350;
        test_data[2595] = 33'd7402090805;
        test_addr[2596] = 351;
        test_data[2596] = 33'd3124014635;
        test_addr[2597] = 352;
        test_data[2597] = 33'd3547444809;
        test_addr[2598] = 353;
        test_data[2598] = 33'd6462933766;
        test_addr[2599] = 354;
        test_data[2599] = 33'd701425537;
        test_addr[2600] = 355;
        test_data[2600] = 33'd1464179666;
        test_addr[2601] = 356;
        test_data[2601] = 33'd2020066253;
        test_addr[2602] = 357;
        test_data[2602] = 33'd2689443698;
        test_addr[2603] = 358;
        test_data[2603] = 33'd2161533557;
        test_addr[2604] = 359;
        test_data[2604] = 33'd4305857401;
        test_addr[2605] = 360;
        test_data[2605] = 33'd1452465810;
        test_addr[2606] = 361;
        test_data[2606] = 33'd3996408431;
        test_addr[2607] = 362;
        test_data[2607] = 33'd2841382309;
        test_addr[2608] = 363;
        test_data[2608] = 33'd2860804675;
        test_addr[2609] = 364;
        test_data[2609] = 33'd1806000219;
        test_addr[2610] = 365;
        test_data[2610] = 33'd3327965930;
        test_addr[2611] = 366;
        test_data[2611] = 33'd3707227066;
        test_addr[2612] = 367;
        test_data[2612] = 33'd1471019555;
        test_addr[2613] = 368;
        test_data[2613] = 33'd1904378792;
        test_addr[2614] = 369;
        test_data[2614] = 33'd2915294719;
        test_addr[2615] = 35;
        test_data[2615] = 33'd5365334139;
        test_addr[2616] = 36;
        test_data[2616] = 33'd946853901;
        test_addr[2617] = 37;
        test_data[2617] = 33'd2604962179;
        test_addr[2618] = 38;
        test_data[2618] = 33'd300770812;
        test_addr[2619] = 39;
        test_data[2619] = 33'd1894311650;
        test_addr[2620] = 40;
        test_data[2620] = 33'd651251042;
        test_addr[2621] = 41;
        test_data[2621] = 33'd3582516170;
        test_addr[2622] = 42;
        test_data[2622] = 33'd2637668923;
        test_addr[2623] = 370;
        test_data[2623] = 33'd1041307001;
        test_addr[2624] = 301;
        test_data[2624] = 33'd2660948838;
        test_addr[2625] = 302;
        test_data[2625] = 33'd2718330062;
        test_addr[2626] = 303;
        test_data[2626] = 33'd1665577570;
        test_addr[2627] = 304;
        test_data[2627] = 33'd3546260524;
        test_addr[2628] = 305;
        test_data[2628] = 33'd409346136;
        test_addr[2629] = 306;
        test_data[2629] = 33'd621355406;
        test_addr[2630] = 307;
        test_data[2630] = 33'd299096324;
        test_addr[2631] = 308;
        test_data[2631] = 33'd3983220710;
        test_addr[2632] = 309;
        test_data[2632] = 33'd4696328025;
        test_addr[2633] = 310;
        test_data[2633] = 33'd6038094765;
        test_addr[2634] = 311;
        test_data[2634] = 33'd3158301700;
        test_addr[2635] = 312;
        test_data[2635] = 33'd3915746261;
        test_addr[2636] = 313;
        test_data[2636] = 33'd494624070;
        test_addr[2637] = 314;
        test_data[2637] = 33'd4281887284;
        test_addr[2638] = 315;
        test_data[2638] = 33'd1927171388;
        test_addr[2639] = 316;
        test_data[2639] = 33'd2860683439;
        test_addr[2640] = 317;
        test_data[2640] = 33'd566819812;
        test_addr[2641] = 318;
        test_data[2641] = 33'd3655450011;
        test_addr[2642] = 319;
        test_data[2642] = 33'd8531489422;
        test_addr[2643] = 320;
        test_data[2643] = 33'd1900882518;
        test_addr[2644] = 321;
        test_data[2644] = 33'd1570807058;
        test_addr[2645] = 322;
        test_data[2645] = 33'd6741247693;
        test_addr[2646] = 323;
        test_data[2646] = 33'd5844198302;
        test_addr[2647] = 324;
        test_data[2647] = 33'd1485894970;
        test_addr[2648] = 325;
        test_data[2648] = 33'd8152587405;
        test_addr[2649] = 326;
        test_data[2649] = 33'd7617320684;
        test_addr[2650] = 327;
        test_data[2650] = 33'd3743832391;
        test_addr[2651] = 328;
        test_data[2651] = 33'd7556934820;
        test_addr[2652] = 329;
        test_data[2652] = 33'd4274943931;
        test_addr[2653] = 330;
        test_data[2653] = 33'd1201882390;
        test_addr[2654] = 331;
        test_data[2654] = 33'd438139954;
        test_addr[2655] = 332;
        test_data[2655] = 33'd1967670189;
        test_addr[2656] = 333;
        test_data[2656] = 33'd1019459317;
        test_addr[2657] = 334;
        test_data[2657] = 33'd1631873129;
        test_addr[2658] = 335;
        test_data[2658] = 33'd1584041641;
        test_addr[2659] = 336;
        test_data[2659] = 33'd5061823108;
        test_addr[2660] = 337;
        test_data[2660] = 33'd5826776752;
        test_addr[2661] = 371;
        test_data[2661] = 33'd7686931035;
        test_addr[2662] = 372;
        test_data[2662] = 33'd2201148884;
        test_addr[2663] = 373;
        test_data[2663] = 33'd7839853763;
        test_addr[2664] = 374;
        test_data[2664] = 33'd86209782;
        test_addr[2665] = 375;
        test_data[2665] = 33'd1901980509;
        test_addr[2666] = 376;
        test_data[2666] = 33'd7217254326;
        test_addr[2667] = 377;
        test_data[2667] = 33'd7885824105;
        test_addr[2668] = 338;
        test_data[2668] = 33'd8214067399;
        test_addr[2669] = 378;
        test_data[2669] = 33'd1303994115;
        test_addr[2670] = 379;
        test_data[2670] = 33'd3489286605;
        test_addr[2671] = 380;
        test_data[2671] = 33'd909919624;
        test_addr[2672] = 65;
        test_data[2672] = 33'd1242253442;
        test_addr[2673] = 381;
        test_data[2673] = 33'd7258224833;
        test_addr[2674] = 382;
        test_data[2674] = 33'd2070296687;
        test_addr[2675] = 383;
        test_data[2675] = 33'd4332516052;
        test_addr[2676] = 384;
        test_data[2676] = 33'd1787421458;
        test_addr[2677] = 385;
        test_data[2677] = 33'd7798665256;
        test_addr[2678] = 386;
        test_data[2678] = 33'd1757687415;
        test_addr[2679] = 387;
        test_data[2679] = 33'd6724848161;
        test_addr[2680] = 388;
        test_data[2680] = 33'd2794749959;
        test_addr[2681] = 389;
        test_data[2681] = 33'd3611635867;
        test_addr[2682] = 390;
        test_data[2682] = 33'd1980103462;
        test_addr[2683] = 391;
        test_data[2683] = 33'd2712963902;
        test_addr[2684] = 392;
        test_data[2684] = 33'd1088256129;
        test_addr[2685] = 393;
        test_data[2685] = 33'd7504250982;
        test_addr[2686] = 394;
        test_data[2686] = 33'd862789604;
        test_addr[2687] = 395;
        test_data[2687] = 33'd6910836485;
        test_addr[2688] = 396;
        test_data[2688] = 33'd5658403625;
        test_addr[2689] = 397;
        test_data[2689] = 33'd1575257700;
        test_addr[2690] = 398;
        test_data[2690] = 33'd5366519133;
        test_addr[2691] = 399;
        test_data[2691] = 33'd7862576228;
        test_addr[2692] = 400;
        test_data[2692] = 33'd523664291;
        test_addr[2693] = 401;
        test_data[2693] = 33'd1851728206;
        test_addr[2694] = 402;
        test_data[2694] = 33'd3042682872;
        test_addr[2695] = 403;
        test_data[2695] = 33'd4090748671;
        test_addr[2696] = 791;
        test_data[2696] = 33'd2331669179;
        test_addr[2697] = 792;
        test_data[2697] = 33'd7566939652;
        test_addr[2698] = 793;
        test_data[2698] = 33'd6173869899;
        test_addr[2699] = 794;
        test_data[2699] = 33'd2371798522;
        test_addr[2700] = 795;
        test_data[2700] = 33'd4674381237;
        test_addr[2701] = 796;
        test_data[2701] = 33'd1668815192;
        test_addr[2702] = 797;
        test_data[2702] = 33'd3852826982;
        test_addr[2703] = 798;
        test_data[2703] = 33'd6765493753;
        test_addr[2704] = 799;
        test_data[2704] = 33'd6209078191;
        test_addr[2705] = 800;
        test_data[2705] = 33'd3694851582;
        test_addr[2706] = 801;
        test_data[2706] = 33'd7008530530;
        test_addr[2707] = 802;
        test_data[2707] = 33'd554375062;
        test_addr[2708] = 803;
        test_data[2708] = 33'd2932332547;
        test_addr[2709] = 804;
        test_data[2709] = 33'd3235881523;
        test_addr[2710] = 805;
        test_data[2710] = 33'd6935891575;
        test_addr[2711] = 806;
        test_data[2711] = 33'd3113296974;
        test_addr[2712] = 807;
        test_data[2712] = 33'd1709814211;
        test_addr[2713] = 808;
        test_data[2713] = 33'd3076343433;
        test_addr[2714] = 809;
        test_data[2714] = 33'd31195618;
        test_addr[2715] = 810;
        test_data[2715] = 33'd1184144647;
        test_addr[2716] = 811;
        test_data[2716] = 33'd3621820777;
        test_addr[2717] = 812;
        test_data[2717] = 33'd2940558418;
        test_addr[2718] = 813;
        test_data[2718] = 33'd5012473762;
        test_addr[2719] = 814;
        test_data[2719] = 33'd6985660589;
        test_addr[2720] = 815;
        test_data[2720] = 33'd7472277175;
        test_addr[2721] = 816;
        test_data[2721] = 33'd96275483;
        test_addr[2722] = 817;
        test_data[2722] = 33'd1666061305;
        test_addr[2723] = 818;
        test_data[2723] = 33'd6375030826;
        test_addr[2724] = 819;
        test_data[2724] = 33'd1667358040;
        test_addr[2725] = 820;
        test_data[2725] = 33'd3676412073;
        test_addr[2726] = 821;
        test_data[2726] = 33'd707615435;
        test_addr[2727] = 822;
        test_data[2727] = 33'd2246158781;
        test_addr[2728] = 823;
        test_data[2728] = 33'd3638573662;
        test_addr[2729] = 824;
        test_data[2729] = 33'd2978602516;
        test_addr[2730] = 825;
        test_data[2730] = 33'd276834200;
        test_addr[2731] = 826;
        test_data[2731] = 33'd1588366455;
        test_addr[2732] = 827;
        test_data[2732] = 33'd481387705;
        test_addr[2733] = 828;
        test_data[2733] = 33'd4327974483;
        test_addr[2734] = 829;
        test_data[2734] = 33'd7115142369;
        test_addr[2735] = 830;
        test_data[2735] = 33'd2929608453;
        test_addr[2736] = 404;
        test_data[2736] = 33'd478746838;
        test_addr[2737] = 405;
        test_data[2737] = 33'd8542882242;
        test_addr[2738] = 406;
        test_data[2738] = 33'd2076323601;
        test_addr[2739] = 407;
        test_data[2739] = 33'd7757891783;
        test_addr[2740] = 547;
        test_data[2740] = 33'd4947557382;
        test_addr[2741] = 548;
        test_data[2741] = 33'd3807612461;
        test_addr[2742] = 549;
        test_data[2742] = 33'd2484022925;
        test_addr[2743] = 550;
        test_data[2743] = 33'd2131016181;
        test_addr[2744] = 551;
        test_data[2744] = 33'd4294945315;
        test_addr[2745] = 552;
        test_data[2745] = 33'd3583226745;
        test_addr[2746] = 553;
        test_data[2746] = 33'd4496330490;
        test_addr[2747] = 408;
        test_data[2747] = 33'd4272217241;
        test_addr[2748] = 409;
        test_data[2748] = 33'd2962982112;
        test_addr[2749] = 410;
        test_data[2749] = 33'd327705331;
        test_addr[2750] = 411;
        test_data[2750] = 33'd1638656261;
        test_addr[2751] = 412;
        test_data[2751] = 33'd1831501086;
        test_addr[2752] = 413;
        test_data[2752] = 33'd3893899942;
        test_addr[2753] = 414;
        test_data[2753] = 33'd1927908942;
        test_addr[2754] = 415;
        test_data[2754] = 33'd3159116717;
        test_addr[2755] = 416;
        test_data[2755] = 33'd1219202730;
        test_addr[2756] = 417;
        test_data[2756] = 33'd2011382593;
        test_addr[2757] = 472;
        test_data[2757] = 33'd7386127003;
        test_addr[2758] = 473;
        test_data[2758] = 33'd6924333958;
        test_addr[2759] = 474;
        test_data[2759] = 33'd8293922366;
        test_addr[2760] = 475;
        test_data[2760] = 33'd3259448472;
        test_addr[2761] = 476;
        test_data[2761] = 33'd3314836530;
        test_addr[2762] = 477;
        test_data[2762] = 33'd4810702126;
        test_addr[2763] = 418;
        test_data[2763] = 33'd5954735385;
        test_addr[2764] = 419;
        test_data[2764] = 33'd3199330442;
        test_addr[2765] = 420;
        test_data[2765] = 33'd6290095488;
        test_addr[2766] = 421;
        test_data[2766] = 33'd1376576240;
        test_addr[2767] = 422;
        test_data[2767] = 33'd712524200;
        test_addr[2768] = 423;
        test_data[2768] = 33'd7591750489;
        test_addr[2769] = 548;
        test_data[2769] = 33'd7287626027;
        test_addr[2770] = 549;
        test_data[2770] = 33'd2484022925;
        test_addr[2771] = 550;
        test_data[2771] = 33'd2131016181;
        test_addr[2772] = 551;
        test_data[2772] = 33'd6951983952;
        test_addr[2773] = 552;
        test_data[2773] = 33'd7563289508;
        test_addr[2774] = 553;
        test_data[2774] = 33'd5231404270;
        test_addr[2775] = 554;
        test_data[2775] = 33'd7445780030;
        test_addr[2776] = 555;
        test_data[2776] = 33'd4696542552;
        test_addr[2777] = 556;
        test_data[2777] = 33'd174607435;
        test_addr[2778] = 424;
        test_data[2778] = 33'd5654680455;
        test_addr[2779] = 425;
        test_data[2779] = 33'd4239458745;
        test_addr[2780] = 426;
        test_data[2780] = 33'd4531632087;
        test_addr[2781] = 427;
        test_data[2781] = 33'd2317805874;
        test_addr[2782] = 428;
        test_data[2782] = 33'd3161887892;
        test_addr[2783] = 429;
        test_data[2783] = 33'd523036013;
        test_addr[2784] = 430;
        test_data[2784] = 33'd4102642570;
        test_addr[2785] = 431;
        test_data[2785] = 33'd245955697;
        test_addr[2786] = 432;
        test_data[2786] = 33'd4738179635;
        test_addr[2787] = 433;
        test_data[2787] = 33'd8355799982;
        test_addr[2788] = 434;
        test_data[2788] = 33'd4623133480;
        test_addr[2789] = 435;
        test_data[2789] = 33'd6749190241;
        test_addr[2790] = 436;
        test_data[2790] = 33'd6420256619;
        test_addr[2791] = 437;
        test_data[2791] = 33'd2623801413;
        test_addr[2792] = 920;
        test_data[2792] = 33'd3297248776;
        test_addr[2793] = 921;
        test_data[2793] = 33'd7572719733;
        test_addr[2794] = 922;
        test_data[2794] = 33'd268862713;
        test_addr[2795] = 923;
        test_data[2795] = 33'd2554414221;
        test_addr[2796] = 924;
        test_data[2796] = 33'd6405337198;
        test_addr[2797] = 925;
        test_data[2797] = 33'd4463869414;
        test_addr[2798] = 438;
        test_data[2798] = 33'd5868618273;
        test_addr[2799] = 439;
        test_data[2799] = 33'd4263494862;
        test_addr[2800] = 440;
        test_data[2800] = 33'd5855248712;
        test_addr[2801] = 441;
        test_data[2801] = 33'd6689078201;
        test_addr[2802] = 442;
        test_data[2802] = 33'd1182124915;
        test_addr[2803] = 443;
        test_data[2803] = 33'd5559814391;
        test_addr[2804] = 444;
        test_data[2804] = 33'd4955300400;
        test_addr[2805] = 445;
        test_data[2805] = 33'd4020894215;
        test_addr[2806] = 578;
        test_data[2806] = 33'd741309116;
        test_addr[2807] = 579;
        test_data[2807] = 33'd3286825499;
        test_addr[2808] = 580;
        test_data[2808] = 33'd376561783;
        test_addr[2809] = 581;
        test_data[2809] = 33'd5597897246;
        test_addr[2810] = 582;
        test_data[2810] = 33'd6515642127;
        test_addr[2811] = 583;
        test_data[2811] = 33'd6816973135;
        test_addr[2812] = 584;
        test_data[2812] = 33'd6226279684;
        test_addr[2813] = 585;
        test_data[2813] = 33'd1415357636;
        test_addr[2814] = 586;
        test_data[2814] = 33'd3407577517;
        test_addr[2815] = 587;
        test_data[2815] = 33'd5250941045;
        test_addr[2816] = 588;
        test_data[2816] = 33'd1568993292;
        test_addr[2817] = 589;
        test_data[2817] = 33'd2295885502;
        test_addr[2818] = 590;
        test_data[2818] = 33'd7337172916;
        test_addr[2819] = 591;
        test_data[2819] = 33'd720614045;
        test_addr[2820] = 592;
        test_data[2820] = 33'd667391101;
        test_addr[2821] = 593;
        test_data[2821] = 33'd3272624999;
        test_addr[2822] = 594;
        test_data[2822] = 33'd5218360596;
        test_addr[2823] = 595;
        test_data[2823] = 33'd6456016398;
        test_addr[2824] = 596;
        test_data[2824] = 33'd7358177755;
        test_addr[2825] = 597;
        test_data[2825] = 33'd6415299630;
        test_addr[2826] = 598;
        test_data[2826] = 33'd7768394115;
        test_addr[2827] = 599;
        test_data[2827] = 33'd3752407160;
        test_addr[2828] = 600;
        test_data[2828] = 33'd3556822102;
        test_addr[2829] = 601;
        test_data[2829] = 33'd6535872974;
        test_addr[2830] = 602;
        test_data[2830] = 33'd996691828;
        test_addr[2831] = 603;
        test_data[2831] = 33'd8177461050;
        test_addr[2832] = 604;
        test_data[2832] = 33'd7284407175;
        test_addr[2833] = 605;
        test_data[2833] = 33'd4062492645;
        test_addr[2834] = 606;
        test_data[2834] = 33'd5957150897;
        test_addr[2835] = 607;
        test_data[2835] = 33'd2708199527;
        test_addr[2836] = 608;
        test_data[2836] = 33'd670098572;
        test_addr[2837] = 609;
        test_data[2837] = 33'd412456713;
        test_addr[2838] = 610;
        test_data[2838] = 33'd3240265434;
        test_addr[2839] = 446;
        test_data[2839] = 33'd2862511605;
        test_addr[2840] = 447;
        test_data[2840] = 33'd5036202736;
        test_addr[2841] = 448;
        test_data[2841] = 33'd7983856578;
        test_addr[2842] = 449;
        test_data[2842] = 33'd3800756962;
        test_addr[2843] = 450;
        test_data[2843] = 33'd3977574422;
        test_addr[2844] = 451;
        test_data[2844] = 33'd8035679255;
        test_addr[2845] = 452;
        test_data[2845] = 33'd343985587;
        test_addr[2846] = 453;
        test_data[2846] = 33'd5216013790;
        test_addr[2847] = 454;
        test_data[2847] = 33'd3300158188;
        test_addr[2848] = 455;
        test_data[2848] = 33'd6605317055;
        test_addr[2849] = 456;
        test_data[2849] = 33'd5635013827;
        test_addr[2850] = 457;
        test_data[2850] = 33'd6456284193;
        test_addr[2851] = 599;
        test_data[2851] = 33'd5179379971;
        test_addr[2852] = 600;
        test_data[2852] = 33'd3556822102;
        test_addr[2853] = 601;
        test_data[2853] = 33'd2240905678;
        test_addr[2854] = 602;
        test_data[2854] = 33'd996691828;
        test_addr[2855] = 603;
        test_data[2855] = 33'd8048775100;
        test_addr[2856] = 604;
        test_data[2856] = 33'd2989439879;
        test_addr[2857] = 605;
        test_data[2857] = 33'd5505638036;
        test_addr[2858] = 606;
        test_data[2858] = 33'd1662183601;
        test_addr[2859] = 607;
        test_data[2859] = 33'd2708199527;
        test_addr[2860] = 458;
        test_data[2860] = 33'd903983808;
        test_addr[2861] = 459;
        test_data[2861] = 33'd600779198;
        test_addr[2862] = 460;
        test_data[2862] = 33'd2637259332;
        test_addr[2863] = 461;
        test_data[2863] = 33'd463249756;
        test_addr[2864] = 462;
        test_data[2864] = 33'd1387176348;
        test_addr[2865] = 463;
        test_data[2865] = 33'd4096796069;
        test_addr[2866] = 464;
        test_data[2866] = 33'd4963550311;
        test_addr[2867] = 465;
        test_data[2867] = 33'd2637855582;
        test_addr[2868] = 1005;
        test_data[2868] = 33'd800335797;
        test_addr[2869] = 1006;
        test_data[2869] = 33'd6115810224;
        test_addr[2870] = 1007;
        test_data[2870] = 33'd492031920;
        test_addr[2871] = 1008;
        test_data[2871] = 33'd2946475741;
        test_addr[2872] = 1009;
        test_data[2872] = 33'd5562244051;
        test_addr[2873] = 1010;
        test_data[2873] = 33'd7608677227;
        test_addr[2874] = 1011;
        test_data[2874] = 33'd1029461814;
        test_addr[2875] = 1012;
        test_data[2875] = 33'd3692205187;
        test_addr[2876] = 1013;
        test_data[2876] = 33'd2547033048;
        test_addr[2877] = 1014;
        test_data[2877] = 33'd1358387716;
        test_addr[2878] = 1015;
        test_data[2878] = 33'd2574971247;
        test_addr[2879] = 1016;
        test_data[2879] = 33'd5401477053;
        test_addr[2880] = 1017;
        test_data[2880] = 33'd4080120458;
        test_addr[2881] = 1018;
        test_data[2881] = 33'd6159364184;
        test_addr[2882] = 1019;
        test_data[2882] = 33'd7922481296;
        test_addr[2883] = 1020;
        test_data[2883] = 33'd6665882113;
        test_addr[2884] = 1021;
        test_data[2884] = 33'd23045195;
        test_addr[2885] = 1022;
        test_data[2885] = 33'd1277705246;
        test_addr[2886] = 1023;
        test_data[2886] = 33'd2086004592;
        test_addr[2887] = 0;
        test_data[2887] = 33'd812361294;
        test_addr[2888] = 1;
        test_data[2888] = 33'd1897396466;
        test_addr[2889] = 2;
        test_data[2889] = 33'd1865453439;
        test_addr[2890] = 3;
        test_data[2890] = 33'd7685124086;
        test_addr[2891] = 4;
        test_data[2891] = 33'd93557296;
        test_addr[2892] = 5;
        test_data[2892] = 33'd838687445;
        test_addr[2893] = 6;
        test_data[2893] = 33'd7690789556;
        test_addr[2894] = 7;
        test_data[2894] = 33'd6853405312;
        test_addr[2895] = 8;
        test_data[2895] = 33'd6568299978;
        test_addr[2896] = 9;
        test_data[2896] = 33'd4367992616;
        test_addr[2897] = 10;
        test_data[2897] = 33'd1664182063;
        test_addr[2898] = 11;
        test_data[2898] = 33'd4491075259;
        test_addr[2899] = 12;
        test_data[2899] = 33'd3296343955;
        test_addr[2900] = 13;
        test_data[2900] = 33'd4630404432;
        test_addr[2901] = 466;
        test_data[2901] = 33'd6838439876;
        test_addr[2902] = 467;
        test_data[2902] = 33'd579888698;
        test_addr[2903] = 468;
        test_data[2903] = 33'd229599703;
        test_addr[2904] = 469;
        test_data[2904] = 33'd3916533083;
        test_addr[2905] = 470;
        test_data[2905] = 33'd3758623902;
        test_addr[2906] = 471;
        test_data[2906] = 33'd4277788026;
        test_addr[2907] = 472;
        test_data[2907] = 33'd3091159707;
        test_addr[2908] = 473;
        test_data[2908] = 33'd7524820018;
        test_addr[2909] = 474;
        test_data[2909] = 33'd3998955070;
        test_addr[2910] = 475;
        test_data[2910] = 33'd7238330659;
        test_addr[2911] = 625;
        test_data[2911] = 33'd6850758234;
        test_addr[2912] = 626;
        test_data[2912] = 33'd3713789991;
        test_addr[2913] = 627;
        test_data[2913] = 33'd8356005006;
        test_addr[2914] = 628;
        test_data[2914] = 33'd3449788833;
        test_addr[2915] = 629;
        test_data[2915] = 33'd1317727169;
        test_addr[2916] = 630;
        test_data[2916] = 33'd3548473177;
        test_addr[2917] = 631;
        test_data[2917] = 33'd7508290992;
        test_addr[2918] = 632;
        test_data[2918] = 33'd173501673;
        test_addr[2919] = 633;
        test_data[2919] = 33'd2419434228;
        test_addr[2920] = 634;
        test_data[2920] = 33'd5158345414;
        test_addr[2921] = 635;
        test_data[2921] = 33'd8443145434;
        test_addr[2922] = 476;
        test_data[2922] = 33'd3314836530;
        test_addr[2923] = 477;
        test_data[2923] = 33'd515734830;
        test_addr[2924] = 478;
        test_data[2924] = 33'd3938658140;
        test_addr[2925] = 479;
        test_data[2925] = 33'd6691164899;
        test_addr[2926] = 480;
        test_data[2926] = 33'd6212319975;
        test_addr[2927] = 481;
        test_data[2927] = 33'd3956236381;
        test_addr[2928] = 482;
        test_data[2928] = 33'd3069633443;
        test_addr[2929] = 483;
        test_data[2929] = 33'd2649187208;
        test_addr[2930] = 484;
        test_data[2930] = 33'd4269737784;
        test_addr[2931] = 485;
        test_data[2931] = 33'd3345226134;
        test_addr[2932] = 486;
        test_data[2932] = 33'd1324217527;
        test_addr[2933] = 487;
        test_data[2933] = 33'd6774294850;
        test_addr[2934] = 488;
        test_data[2934] = 33'd5358175234;
        test_addr[2935] = 489;
        test_data[2935] = 33'd3950820746;
        test_addr[2936] = 490;
        test_data[2936] = 33'd3214783106;
        test_addr[2937] = 491;
        test_data[2937] = 33'd7279381255;
        test_addr[2938] = 492;
        test_data[2938] = 33'd1809665157;
        test_addr[2939] = 493;
        test_data[2939] = 33'd879737958;
        test_addr[2940] = 494;
        test_data[2940] = 33'd821347042;
        test_addr[2941] = 495;
        test_data[2941] = 33'd7613236433;
        test_addr[2942] = 496;
        test_data[2942] = 33'd3581785694;
        test_addr[2943] = 497;
        test_data[2943] = 33'd1177368502;
        test_addr[2944] = 498;
        test_data[2944] = 33'd3822144455;
        test_addr[2945] = 499;
        test_data[2945] = 33'd3997100319;
        test_addr[2946] = 500;
        test_data[2946] = 33'd6491033823;
        test_addr[2947] = 501;
        test_data[2947] = 33'd6507984027;
        test_addr[2948] = 502;
        test_data[2948] = 33'd1457378795;
        test_addr[2949] = 503;
        test_data[2949] = 33'd13805880;
        test_addr[2950] = 504;
        test_data[2950] = 33'd2586581290;
        test_addr[2951] = 505;
        test_data[2951] = 33'd7339973833;
        test_addr[2952] = 154;
        test_data[2952] = 33'd6864757999;
        test_addr[2953] = 506;
        test_data[2953] = 33'd2189946085;
        test_addr[2954] = 507;
        test_data[2954] = 33'd790225939;
        test_addr[2955] = 508;
        test_data[2955] = 33'd750930004;
        test_addr[2956] = 509;
        test_data[2956] = 33'd4443750001;
        test_addr[2957] = 510;
        test_data[2957] = 33'd1738761925;
        test_addr[2958] = 511;
        test_data[2958] = 33'd868517225;
        test_addr[2959] = 512;
        test_data[2959] = 33'd3634725493;
        test_addr[2960] = 513;
        test_data[2960] = 33'd45075662;
        test_addr[2961] = 514;
        test_data[2961] = 33'd3808305303;
        test_addr[2962] = 515;
        test_data[2962] = 33'd934899158;
        test_addr[2963] = 516;
        test_data[2963] = 33'd3277394190;
        test_addr[2964] = 438;
        test_data[2964] = 33'd1573650977;
        test_addr[2965] = 439;
        test_data[2965] = 33'd7753752820;
        test_addr[2966] = 440;
        test_data[2966] = 33'd1560281416;
        test_addr[2967] = 441;
        test_data[2967] = 33'd5826272205;
        test_addr[2968] = 442;
        test_data[2968] = 33'd7112344951;
        test_addr[2969] = 443;
        test_data[2969] = 33'd5915776467;
        test_addr[2970] = 444;
        test_data[2970] = 33'd660333104;
        test_addr[2971] = 445;
        test_data[2971] = 33'd4020894215;
        test_addr[2972] = 446;
        test_data[2972] = 33'd2862511605;
        test_addr[2973] = 447;
        test_data[2973] = 33'd741235440;
        test_addr[2974] = 448;
        test_data[2974] = 33'd8302971071;
        test_addr[2975] = 517;
        test_data[2975] = 33'd8317199872;
        test_addr[2976] = 518;
        test_data[2976] = 33'd209533787;
        test_addr[2977] = 519;
        test_data[2977] = 33'd5747125812;
        test_addr[2978] = 520;
        test_data[2978] = 33'd4515879748;
        test_addr[2979] = 238;
        test_data[2979] = 33'd736219013;
        test_addr[2980] = 239;
        test_data[2980] = 33'd1052350388;
        test_addr[2981] = 240;
        test_data[2981] = 33'd7132222017;
        test_addr[2982] = 241;
        test_data[2982] = 33'd8139133701;
        test_addr[2983] = 242;
        test_data[2983] = 33'd2915968114;
        test_addr[2984] = 243;
        test_data[2984] = 33'd6032243847;
        test_addr[2985] = 521;
        test_data[2985] = 33'd1168067242;
        test_addr[2986] = 522;
        test_data[2986] = 33'd6509343582;
        test_addr[2987] = 523;
        test_data[2987] = 33'd5101737760;
        test_addr[2988] = 524;
        test_data[2988] = 33'd3720168166;
        test_addr[2989] = 525;
        test_data[2989] = 33'd2968836141;
        test_addr[2990] = 526;
        test_data[2990] = 33'd2513327218;
        test_addr[2991] = 527;
        test_data[2991] = 33'd7141611420;
        test_addr[2992] = 528;
        test_data[2992] = 33'd7776663827;
        test_addr[2993] = 529;
        test_data[2993] = 33'd3177420342;
        test_addr[2994] = 530;
        test_data[2994] = 33'd677310380;
        test_addr[2995] = 531;
        test_data[2995] = 33'd4269338406;
        test_addr[2996] = 532;
        test_data[2996] = 33'd1758387349;
        test_addr[2997] = 533;
        test_data[2997] = 33'd4804837348;
        test_addr[2998] = 534;
        test_data[2998] = 33'd6923391952;
        test_addr[2999] = 535;
        test_data[2999] = 33'd7196258704;

    end
endmodule


`timescale 1ns/1ps
module mem_bram #(
    parameter ADDR_WIDTH = 10,		//地址宽度
    parameter DATA_WIDTH = 128		//数据宽度
)(
    input                   clk,   // Clock
    input [ADDR_WIDTH-1:0]  raddr,  // Address
    input [ADDR_WIDTH-1:0]  waddr,  // Address
    input [DATA_WIDTH-1:0]  din,   // Data Input
    input                   we,    // Write Enable
    output [DATA_WIDTH-1:0] dout   // Data Output
); 
    reg [ADDR_WIDTH-1:0] addr_r;  // Address Register
    reg [DATA_WIDTH-1:0] ram [0:(1 << ADDR_WIDTH)-1];
    integer i;
    initial begin
        ram[0][31:0] = 32'd812361294;
        ram[0][63:32] = 32'd1897396466;
        ram[0][95:64] = 32'd3157995732;
        ram[0][127:96] = 32'd3965266920;
        ram[1][31:0] = 32'd164470890;
        ram[1][63:32] = 32'd4813263;
        ram[1][95:64] = 32'd1309544095;
        ram[1][127:96] = 32'd3491080214;
        ram[2][31:0] = 32'd1793239769;
        ram[2][63:32] = 32'd1174159001;
        ram[2][95:64] = 32'd1664182063;
        ram[2][127:96] = 32'd773081521;
        ram[3][31:0] = 32'd3296343955;
        ram[3][63:32] = 32'd1476987912;
        ram[3][95:64] = 32'd1747019271;
        ram[3][127:96] = 32'd2749577582;
        ram[4][31:0] = 32'd2962149009;
        ram[4][63:32] = 32'd1707974702;
        ram[4][95:64] = 32'd2033398483;
        ram[4][127:96] = 32'd1943724055;
        ram[5][31:0] = 32'd1223440380;
        ram[5][63:32] = 32'd3366782182;
        ram[5][95:64] = 32'd883716006;
        ram[5][127:96] = 32'd2361297799;
        ram[6][31:0] = 32'd2711593210;
        ram[6][63:32] = 32'd4002336428;
        ram[6][95:64] = 32'd4291600053;
        ram[6][127:96] = 32'd4190492404;
        ram[7][31:0] = 32'd1899814066;
        ram[7][63:32] = 32'd3331445440;
        ram[7][95:64] = 32'd1741498846;
        ram[7][127:96] = 32'd3230234606;
        ram[8][31:0] = 32'd1170076186;
        ram[8][63:32] = 32'd2359621732;
        ram[8][95:64] = 32'd1887051034;
        ram[8][127:96] = 32'd2113332559;
        ram[9][31:0] = 32'd2709550290;
        ram[9][63:32] = 32'd406326701;
        ram[9][95:64] = 32'd3133901872;
        ram[9][127:96] = 32'd1715945728;
        ram[10][31:0] = 32'd3642725099;
        ram[10][63:32] = 32'd2411058451;
        ram[10][95:64] = 32'd3969759003;
        ram[10][127:96] = 32'd389770497;
        ram[11][31:0] = 32'd2890247156;
        ram[11][63:32] = 32'd1444532856;
        ram[11][95:64] = 32'd2921447489;
        ram[11][127:96] = 32'd3675966926;
        ram[12][31:0] = 32'd64235302;
        ram[12][63:32] = 32'd1390656163;
        ram[12][95:64] = 32'd2480296893;
        ram[12][127:96] = 32'd893530107;
        ram[13][31:0] = 32'd369651485;
        ram[13][63:32] = 32'd2187729913;
        ram[13][95:64] = 32'd1681690332;
        ram[13][127:96] = 32'd1478733057;
        ram[14][31:0] = 32'd13033719;
        ram[14][63:32] = 32'd691835738;
        ram[14][95:64] = 32'd528146972;
        ram[14][127:96] = 32'd106529920;
        ram[15][31:0] = 32'd2587167315;
        ram[15][63:32] = 32'd3444518270;
        ram[15][95:64] = 32'd2627318154;
        ram[15][127:96] = 32'd12778738;
        ram[16][31:0] = 32'd4280548596;
        ram[16][63:32] = 32'd3000665519;
        ram[16][95:64] = 32'd2358437066;
        ram[16][127:96] = 32'd1974385293;
        ram[17][31:0] = 32'd1457236560;
        ram[17][63:32] = 32'd912614945;
        ram[17][95:64] = 32'd2389449862;
        ram[17][127:96] = 32'd2460511432;
        ram[18][31:0] = 32'd414705635;
        ram[18][63:32] = 32'd3301388465;
        ram[18][95:64] = 32'd2014563986;
        ram[18][127:96] = 32'd3636478413;
        ram[19][31:0] = 32'd1338201231;
        ram[19][63:32] = 32'd2865448495;
        ram[19][95:64] = 32'd1953052136;
        ram[19][127:96] = 32'd1775955632;
        ram[20][31:0] = 32'd4154877383;
        ram[20][63:32] = 32'd3550050089;
        ram[20][95:64] = 32'd1564001926;
        ram[20][127:96] = 32'd1729932993;
        ram[21][31:0] = 32'd1629692541;
        ram[21][63:32] = 32'd2686387223;
        ram[21][95:64] = 32'd375741016;
        ram[21][127:96] = 32'd405157155;
        ram[22][31:0] = 32'd2879312064;
        ram[22][63:32] = 32'd3559542326;
        ram[22][95:64] = 32'd3551737466;
        ram[22][127:96] = 32'd1285586415;
        ram[23][31:0] = 32'd1656551191;
        ram[23][63:32] = 32'd1856969724;
        ram[23][95:64] = 32'd2987649344;
        ram[23][127:96] = 32'd2737991781;
        ram[24][31:0] = 32'd3739168123;
        ram[24][63:32] = 32'd1649687892;
        ram[24][95:64] = 32'd2397619105;
        ram[24][127:96] = 32'd3659483916;
        ram[25][31:0] = 32'd1882137235;
        ram[25][63:32] = 32'd1616255243;
        ram[25][95:64] = 32'd1662993831;
        ram[25][127:96] = 32'd1019640399;
        ram[26][31:0] = 32'd1424217888;
        ram[26][63:32] = 32'd627517218;
        ram[26][95:64] = 32'd2218451356;
        ram[26][127:96] = 32'd3217439098;
        ram[27][31:0] = 32'd4247265534;
        ram[27][63:32] = 32'd264822472;
        ram[27][95:64] = 32'd4027024129;
        ram[27][127:96] = 32'd645329535;
        ram[28][31:0] = 32'd535433161;
        ram[28][63:32] = 32'd4144529833;
        ram[28][95:64] = 32'd2554819996;
        ram[28][127:96] = 32'd3969435406;
        ram[29][31:0] = 32'd1512917393;
        ram[29][63:32] = 32'd3459749905;
        ram[29][95:64] = 32'd2078089603;
        ram[29][127:96] = 32'd3211090985;
        ram[30][31:0] = 32'd557041591;
        ram[30][63:32] = 32'd3495515776;
        ram[30][95:64] = 32'd886188703;
        ram[30][127:96] = 32'd978523342;
        ram[31][31:0] = 32'd2261534157;
        ram[31][63:32] = 32'd1178766234;
        ram[31][95:64] = 32'd717632510;
        ram[31][127:96] = 32'd2732828399;
        ram[32][31:0] = 32'd1015809205;
        ram[32][63:32] = 32'd438601362;
        ram[32][95:64] = 32'd2760717433;
        ram[32][127:96] = 32'd3219734873;
        ram[33][31:0] = 32'd1457531679;
        ram[33][63:32] = 32'd3756088394;
        ram[33][95:64] = 32'd4205150678;
        ram[33][127:96] = 32'd3470509274;
        ram[34][31:0] = 32'd2230430546;
        ram[34][63:32] = 32'd4277997269;
        ram[34][95:64] = 32'd51940499;
        ram[34][127:96] = 32'd4250352825;
        ram[35][31:0] = 32'd558456538;
        ram[35][63:32] = 32'd485567310;
        ram[35][95:64] = 32'd1458947625;
        ram[35][127:96] = 32'd730436975;
        ram[36][31:0] = 32'd1218308152;
        ram[36][63:32] = 32'd2394330144;
        ram[36][95:64] = 32'd1483917544;
        ram[36][127:96] = 32'd3933851125;
        ram[37][31:0] = 32'd1074274996;
        ram[37][63:32] = 32'd304283732;
        ram[37][95:64] = 32'd1383869392;
        ram[37][127:96] = 32'd2820628440;
        ram[38][31:0] = 32'd112695676;
        ram[38][63:32] = 32'd327985978;
        ram[38][95:64] = 32'd412214464;
        ram[38][127:96] = 32'd3182442945;
        ram[39][31:0] = 32'd4176867573;
        ram[39][63:32] = 32'd1333860272;
        ram[39][95:64] = 32'd4087206092;
        ram[39][127:96] = 32'd4088679797;
        ram[40][31:0] = 32'd347557471;
        ram[40][63:32] = 32'd1498608590;
        ram[40][95:64] = 32'd1461900145;
        ram[40][127:96] = 32'd2045508676;
        ram[41][31:0] = 32'd617221806;
        ram[41][63:32] = 32'd117310100;
        ram[41][95:64] = 32'd2648221725;
        ram[41][127:96] = 32'd142053120;
        ram[42][31:0] = 32'd254554983;
        ram[42][63:32] = 32'd96607098;
        ram[42][95:64] = 32'd574793399;
        ram[42][127:96] = 32'd753209148;
        ram[43][31:0] = 32'd460255681;
        ram[43][63:32] = 32'd4213223392;
        ram[43][95:64] = 32'd1373713971;
        ram[43][127:96] = 32'd1891542300;
        ram[44][31:0] = 32'd2743796502;
        ram[44][63:32] = 32'd1825087556;
        ram[44][95:64] = 32'd3775849174;
        ram[44][127:96] = 32'd1928357839;
        ram[45][31:0] = 32'd3962182398;
        ram[45][63:32] = 32'd1609542177;
        ram[45][95:64] = 32'd557477877;
        ram[45][127:96] = 32'd1320690480;
        ram[46][31:0] = 32'd2515569179;
        ram[46][63:32] = 32'd76388760;
        ram[46][95:64] = 32'd3665623001;
        ram[46][127:96] = 32'd800185981;
        ram[47][31:0] = 32'd3633252065;
        ram[47][63:32] = 32'd3256549792;
        ram[47][95:64] = 32'd3874319877;
        ram[47][127:96] = 32'd4077538423;
        ram[48][31:0] = 32'd1404789710;
        ram[48][63:32] = 32'd2024109334;
        ram[48][95:64] = 32'd117118296;
        ram[48][127:96] = 32'd1198019948;
        ram[49][31:0] = 32'd1622317500;
        ram[49][63:32] = 32'd2750204444;
        ram[49][95:64] = 32'd1532972969;
        ram[49][127:96] = 32'd2378011170;
        ram[50][31:0] = 32'd4250933843;
        ram[50][63:32] = 32'd1833057303;
        ram[50][95:64] = 32'd2638317033;
        ram[50][127:96] = 32'd998547257;
        ram[51][31:0] = 32'd2620591812;
        ram[51][63:32] = 32'd2964469971;
        ram[51][95:64] = 32'd1308783437;
        ram[51][127:96] = 32'd155196010;
        ram[52][31:0] = 32'd1515041615;
        ram[52][63:32] = 32'd3938057574;
        ram[52][95:64] = 32'd2312377961;
        ram[52][127:96] = 32'd2875926310;
        ram[53][31:0] = 32'd2392747211;
        ram[53][63:32] = 32'd3665553539;
        ram[53][95:64] = 32'd1034237452;
        ram[53][127:96] = 32'd2832534662;
        ram[54][31:0] = 32'd2609755010;
        ram[54][63:32] = 32'd1119239002;
        ram[54][95:64] = 32'd2296008684;
        ram[54][127:96] = 32'd3225055293;
        ram[55][31:0] = 32'd1552736584;
        ram[55][63:32] = 32'd1801818893;
        ram[55][95:64] = 32'd727510908;
        ram[55][127:96] = 32'd2764688405;
        ram[56][31:0] = 32'd1983206576;
        ram[56][63:32] = 32'd3019194714;
        ram[56][95:64] = 32'd229751523;
        ram[56][127:96] = 32'd1667423717;
        ram[57][31:0] = 32'd1082603118;
        ram[57][63:32] = 32'd1506219133;
        ram[57][95:64] = 32'd3332009274;
        ram[57][127:96] = 32'd1787072800;
        ram[58][31:0] = 32'd1891418860;
        ram[58][63:32] = 32'd2168623663;
        ram[58][95:64] = 32'd797215018;
        ram[58][127:96] = 32'd3439453128;
        ram[59][31:0] = 32'd795204265;
        ram[59][63:32] = 32'd168920287;
        ram[59][95:64] = 32'd159301787;
        ram[59][127:96] = 32'd3601678559;
        ram[60][31:0] = 32'd3705921312;
        ram[60][63:32] = 32'd1202615656;
        ram[60][95:64] = 32'd1167664452;
        ram[60][127:96] = 32'd874735177;
        ram[61][31:0] = 32'd1146573824;
        ram[61][63:32] = 32'd2038925291;
        ram[61][95:64] = 32'd3389506182;
        ram[61][127:96] = 32'd1086878351;
        ram[62][31:0] = 32'd2433798430;
        ram[62][63:32] = 32'd230942795;
        ram[62][95:64] = 32'd157822933;
        ram[62][127:96] = 32'd2172745435;
        ram[63][31:0] = 32'd3216848485;
        ram[63][63:32] = 32'd522192966;
        ram[63][95:64] = 32'd1000930920;
        ram[63][127:96] = 32'd714439378;
        ram[64][31:0] = 32'd2800244347;
        ram[64][63:32] = 32'd248550902;
        ram[64][95:64] = 32'd3691916876;
        ram[64][127:96] = 32'd2756113887;
        ram[65][31:0] = 32'd1766135903;
        ram[65][63:32] = 32'd4204582623;
        ram[65][95:64] = 32'd1204698417;
        ram[65][127:96] = 32'd2114950029;
        ram[66][31:0] = 32'd823241581;
        ram[66][63:32] = 32'd1728145956;
        ram[66][95:64] = 32'd3223227851;
        ram[66][127:96] = 32'd1691484081;
        ram[67][31:0] = 32'd1602773367;
        ram[67][63:32] = 32'd3034594309;
        ram[67][95:64] = 32'd3716873283;
        ram[67][127:96] = 32'd2102264294;
        ram[68][31:0] = 32'd3539921614;
        ram[68][63:32] = 32'd3701319037;
        ram[68][95:64] = 32'd2004368579;
        ram[68][127:96] = 32'd1824795164;
        ram[69][31:0] = 32'd1921721343;
        ram[69][63:32] = 32'd1860688658;
        ram[69][95:64] = 32'd3515322191;
        ram[69][127:96] = 32'd1883857597;
        ram[70][31:0] = 32'd2299961408;
        ram[70][63:32] = 32'd4110926899;
        ram[70][95:64] = 32'd2071294607;
        ram[70][127:96] = 32'd2622506310;
        ram[71][31:0] = 32'd3230604876;
        ram[71][63:32] = 32'd812304788;
        ram[71][95:64] = 32'd775168527;
        ram[71][127:96] = 32'd2682374959;
        ram[72][31:0] = 32'd1151781196;
        ram[72][63:32] = 32'd2823208990;
        ram[72][95:64] = 32'd2277953385;
        ram[72][127:96] = 32'd1297973981;
        ram[73][31:0] = 32'd273664053;
        ram[73][63:32] = 32'd688835068;
        ram[73][95:64] = 32'd3604100589;
        ram[73][127:96] = 32'd2347942712;
        ram[74][31:0] = 32'd1233127960;
        ram[74][63:32] = 32'd3955483560;
        ram[74][95:64] = 32'd703519346;
        ram[74][127:96] = 32'd3010600461;
        ram[75][31:0] = 32'd1320963640;
        ram[75][63:32] = 32'd2660948838;
        ram[75][95:64] = 32'd1512656212;
        ram[75][127:96] = 32'd3928629502;
        ram[76][31:0] = 32'd861935821;
        ram[76][63:32] = 32'd2556845885;
        ram[76][95:64] = 32'd621355406;
        ram[76][127:96] = 32'd2335768031;
        ram[77][31:0] = 32'd3983220710;
        ram[77][63:32] = 32'd3373852337;
        ram[77][95:64] = 32'd3671954381;
        ram[77][127:96] = 32'd2927272024;
        ram[78][31:0] = 32'd3915746261;
        ram[78][63:32] = 32'd494624070;
        ram[78][95:64] = 32'd3309988311;
        ram[78][127:96] = 32'd1132837972;
        ram[79][31:0] = 32'd2910487772;
        ram[79][63:32] = 32'd3066325816;
        ram[79][95:64] = 32'd3655450011;
        ram[79][127:96] = 32'd2771319734;
        ram[80][31:0] = 32'd59000887;
        ram[80][63:32] = 32'd700513712;
        ram[80][95:64] = 32'd223050916;
        ram[80][127:96] = 32'd1549846123;
        ram[81][31:0] = 32'd1485894970;
        ram[81][63:32] = 32'd1503820403;
        ram[81][95:64] = 32'd20706691;
        ram[81][127:96] = 32'd2856799024;
        ram[82][31:0] = 32'd3027590231;
        ram[82][63:32] = 32'd886386958;
        ram[82][95:64] = 32'd1408921763;
        ram[82][127:96] = 32'd1012710083;
        ram[83][31:0] = 32'd3964024451;
        ram[83][63:32] = 32'd2623422963;
        ram[83][95:64] = 32'd1631873129;
        ram[83][127:96] = 32'd3094982513;
        ram[84][31:0] = 32'd604229382;
        ram[84][63:32] = 32'd190701906;
        ram[84][95:64] = 32'd2063414812;
        ram[84][127:96] = 32'd2384267827;
        ram[85][31:0] = 32'd2877406934;
        ram[85][63:32] = 32'd2186863965;
        ram[85][95:64] = 32'd4078357046;
        ram[85][127:96] = 32'd1123238982;
        ram[86][31:0] = 32'd3796226835;
        ram[86][63:32] = 32'd3794021488;
        ram[86][95:64] = 32'd81294826;
        ram[86][127:96] = 32'd1991678289;
        ram[87][31:0] = 32'd926633043;
        ram[87][63:32] = 32'd205161254;
        ram[87][95:64] = 32'd1629934311;
        ram[87][127:96] = 32'd3124014635;
        ram[88][31:0] = 32'd3793842303;
        ram[88][63:32] = 32'd2049664093;
        ram[88][95:64] = 32'd701425537;
        ram[88][127:96] = 32'd2427207363;
        ram[89][31:0] = 32'd2020066253;
        ram[89][63:32] = 32'd2661076722;
        ram[89][95:64] = 32'd2161533557;
        ram[89][127:96] = 32'd2495672481;
        ram[90][31:0] = 32'd1452465810;
        ram[90][63:32] = 32'd3160518389;
        ram[90][95:64] = 32'd2841382309;
        ram[90][127:96] = 32'd3212580707;
        ram[91][31:0] = 32'd2996693876;
        ram[91][63:32] = 32'd152547103;
        ram[91][95:64] = 32'd3707227066;
        ram[91][127:96] = 32'd1471019555;
        ram[92][31:0] = 32'd1294858093;
        ram[92][63:32] = 32'd2915294719;
        ram[92][95:64] = 32'd1041307001;
        ram[92][127:96] = 32'd2929810272;
        ram[93][31:0] = 32'd19502472;
        ram[93][63:32] = 32'd3262680181;
        ram[93][95:64] = 32'd86209782;
        ram[93][127:96] = 32'd3820989693;
        ram[94][31:0] = 32'd2739596899;
        ram[94][63:32] = 32'd528252277;
        ram[94][95:64] = 32'd1303994115;
        ram[94][127:96] = 32'd3762588080;
        ram[95][31:0] = 32'd909919624;
        ram[95][63:32] = 32'd2494821825;
        ram[95][95:64] = 32'd2070296687;
        ram[95][127:96] = 32'd489544890;
        ram[96][31:0] = 32'd841967182;
        ram[96][63:32] = 32'd792251059;
        ram[96][95:64] = 32'd1757687415;
        ram[96][127:96] = 32'd3967144044;
        ram[97][31:0] = 32'd2794749959;
        ram[97][63:32] = 32'd3611635867;
        ram[97][95:64] = 32'd1980103462;
        ram[97][127:96] = 32'd4203711356;
        ram[98][31:0] = 32'd1088256129;
        ram[98][63:32] = 32'd2750675278;
        ram[98][95:64] = 32'd862789604;
        ram[98][127:96] = 32'd2126893221;
        ram[99][31:0] = 32'd4286897536;
        ram[99][63:32] = 32'd1575257700;
        ram[99][95:64] = 32'd3564413496;
        ram[99][127:96] = 32'd373361739;
        ram[100][31:0] = 32'd523664291;
        ram[100][63:32] = 32'd486121505;
        ram[100][95:64] = 32'd673171958;
        ram[100][127:96] = 32'd3751867044;
        ram[101][31:0] = 32'd478746838;
        ram[101][63:32] = 32'd2789966675;
        ram[101][95:64] = 32'd272467445;
        ram[101][127:96] = 32'd3655415553;
        ram[102][31:0] = 32'd4272217241;
        ram[102][63:32] = 32'd2962982112;
        ram[102][95:64] = 32'd327705331;
        ram[102][127:96] = 32'd1638656261;
        ram[103][31:0] = 32'd1831501086;
        ram[103][63:32] = 32'd3893899942;
        ram[103][95:64] = 32'd1927908942;
        ram[103][127:96] = 32'd3159116717;
        ram[104][31:0] = 32'd4102174094;
        ram[104][63:32] = 32'd2072738163;
        ram[104][95:64] = 32'd717648603;
        ram[104][127:96] = 32'd2628348997;
        ram[105][31:0] = 32'd2417509630;
        ram[105][63:32] = 32'd1376576240;
        ram[105][95:64] = 32'd712524200;
        ram[105][127:96] = 32'd3658904312;
        ram[106][31:0] = 32'd1503454293;
        ram[106][63:32] = 32'd4239458745;
        ram[106][95:64] = 32'd2181778910;
        ram[106][127:96] = 32'd302461623;
        ram[107][31:0] = 32'd3161887892;
        ram[107][63:32] = 32'd523036013;
        ram[107][95:64] = 32'd4102642570;
        ram[107][127:96] = 32'd3040028192;
        ram[108][31:0] = 32'd1817537658;
        ram[108][63:32] = 32'd131728541;
        ram[108][95:64] = 32'd1334678566;
        ram[108][127:96] = 32'd874658310;
        ram[109][31:0] = 32'd3478059314;
        ram[109][63:32] = 32'd138201149;
        ram[109][95:64] = 32'd2780888181;
        ram[109][127:96] = 32'd4263494862;
        ram[110][31:0] = 32'd3617831507;
        ram[110][63:32] = 32'd4133778867;
        ram[110][95:64] = 32'd1182124915;
        ram[110][127:96] = 32'd887054320;
        ram[111][31:0] = 32'd3362594900;
        ram[111][63:32] = 32'd320890295;
        ram[111][95:64] = 32'd2862511605;
        ram[111][127:96] = 32'd2384680284;
        ram[112][31:0] = 32'd1262035775;
        ram[112][63:32] = 32'd1270840210;
        ram[112][95:64] = 32'd3977574422;
        ram[112][127:96] = 32'd2470246955;
        ram[113][31:0] = 32'd2255354623;
        ram[113][63:32] = 32'd1872832286;
        ram[113][95:64] = 32'd1765327971;
        ram[113][127:96] = 32'd2792297812;
        ram[114][31:0] = 32'd3380440245;
        ram[114][63:32] = 32'd2493892019;
        ram[114][95:64] = 32'd1719765622;
        ram[114][127:96] = 32'd600779198;
        ram[115][31:0] = 32'd2977339794;
        ram[115][63:32] = 32'd1567929911;
        ram[115][95:64] = 32'd1387176348;
        ram[115][127:96] = 32'd4096796069;
        ram[116][31:0] = 32'd1087715771;
        ram[116][63:32] = 32'd2637855582;
        ram[116][95:64] = 32'd2023239053;
        ram[116][127:96] = 32'd579888698;
        ram[117][31:0] = 32'd279675755;
        ram[117][63:32] = 32'd3850513177;
        ram[117][95:64] = 32'd2010324295;
        ram[117][127:96] = 32'd2633924524;
        ram[118][31:0] = 32'd1585350521;
        ram[118][63:32] = 32'd1355422752;
        ram[118][95:64] = 32'd4051137299;
        ram[118][127:96] = 32'd3259448472;
        ram[119][31:0] = 32'd3314836530;
        ram[119][63:32] = 32'd2300423720;
        ram[119][95:64] = 32'd3938658140;
        ram[119][127:96] = 32'd3609861208;
        ram[120][31:0] = 32'd1712226038;
        ram[120][63:32] = 32'd1342983001;
        ram[120][95:64] = 32'd3069633443;
        ram[120][127:96] = 32'd2649187208;
        ram[121][31:0] = 32'd4269737784;
        ram[121][63:32] = 32'd3345226134;
        ram[121][95:64] = 32'd1023397519;
        ram[121][127:96] = 32'd4014581281;
        ram[122][31:0] = 32'd1838682392;
        ram[122][63:32] = 32'd1491360199;
        ram[122][95:64] = 32'd1608490784;
        ram[122][127:96] = 32'd1594847873;
        ram[123][31:0] = 32'd1821644561;
        ram[123][63:32] = 32'd1800880124;
        ram[123][95:64] = 32'd821347042;
        ram[123][127:96] = 32'd2117462048;
        ram[124][31:0] = 32'd3581785694;
        ram[124][63:32] = 32'd1177368502;
        ram[124][95:64] = 32'd3822144455;
        ram[124][127:96] = 32'd3127083966;
        ram[125][31:0] = 32'd100230629;
        ram[125][63:32] = 32'd215543822;
        ram[125][95:64] = 32'd1457378795;
        ram[125][127:96] = 32'd3251093126;
        ram[126][31:0] = 32'd2586581290;
        ram[126][63:32] = 32'd2328699311;
        ram[126][95:64] = 32'd2074859986;
        ram[126][127:96] = 32'd475067250;
        ram[127][31:0] = 32'd3858046342;
        ram[127][63:32] = 32'd2012699169;
        ram[127][95:64] = 32'd1161777028;
        ram[127][127:96] = 32'd868517225;
        ram[128][31:0] = 32'd2330170027;
        ram[128][63:32] = 32'd45075662;
        ram[128][95:64] = 32'd1622445132;
        ram[128][127:96] = 32'd934899158;
        ram[129][31:0] = 32'd157205391;
        ram[129][63:32] = 32'd1106079426;
        ram[129][95:64] = 32'd209533787;
        ram[129][127:96] = 32'd2029500360;
        ram[130][31:0] = 32'd1199393578;
        ram[130][63:32] = 32'd1928735641;
        ram[130][95:64] = 32'd4045583222;
        ram[130][127:96] = 32'd3215894844;
        ram[131][31:0] = 32'd3814837793;
        ram[131][63:32] = 32'd3880037807;
        ram[131][95:64] = 32'd2513327218;
        ram[131][127:96] = 32'd3681101907;
        ram[132][31:0] = 32'd1983832739;
        ram[132][63:32] = 32'd3177420342;
        ram[132][95:64] = 32'd1514028413;
        ram[132][127:96] = 32'd4269338406;
        ram[133][31:0] = 32'd1758387349;
        ram[133][63:32] = 32'd3892039782;
        ram[133][95:64] = 32'd3083492837;
        ram[133][127:96] = 32'd4284361995;
        ram[134][31:0] = 32'd3377477922;
        ram[134][63:32] = 32'd1309125160;
        ram[134][95:64] = 32'd1250172866;
        ram[134][127:96] = 32'd2819209516;
        ram[135][31:0] = 32'd1100314726;
        ram[135][63:32] = 32'd3682747475;
        ram[135][95:64] = 32'd1732119287;
        ram[135][127:96] = 32'd81502868;
        ram[136][31:0] = 32'd2034855529;
        ram[136][63:32] = 32'd3917407985;
        ram[136][95:64] = 32'd2114980159;
        ram[136][127:96] = 32'd3961698218;
        ram[137][31:0] = 32'd3807612461;
        ram[137][63:32] = 32'd2484022925;
        ram[137][95:64] = 32'd2131016181;
        ram[137][127:96] = 32'd4294945315;
        ram[138][31:0] = 32'd3583226745;
        ram[138][63:32] = 32'd81343249;
        ram[138][95:64] = 32'd2981022136;
        ram[138][127:96] = 32'd3198658539;
        ram[139][31:0] = 32'd174607435;
        ram[139][63:32] = 32'd1596273533;
        ram[139][95:64] = 32'd862985215;
        ram[139][127:96] = 32'd2286533469;
        ram[140][31:0] = 32'd2440931925;
        ram[140][63:32] = 32'd2008701872;
        ram[140][95:64] = 32'd1056483800;
        ram[140][127:96] = 32'd1776101444;
        ram[141][31:0] = 32'd2025943392;
        ram[141][63:32] = 32'd3264098589;
        ram[141][95:64] = 32'd1836238996;
        ram[141][127:96] = 32'd2887167439;
        ram[142][31:0] = 32'd2411940668;
        ram[142][63:32] = 32'd2786633091;
        ram[142][95:64] = 32'd3634409579;
        ram[142][127:96] = 32'd2590447935;
        ram[143][31:0] = 32'd3141059683;
        ram[143][63:32] = 32'd4029761842;
        ram[143][95:64] = 32'd4104262188;
        ram[143][127:96] = 32'd197152237;
        ram[144][31:0] = 32'd65320894;
        ram[144][63:32] = 32'd4153629096;
        ram[144][95:64] = 32'd741309116;
        ram[144][127:96] = 32'd1009033767;
        ram[145][31:0] = 32'd3021320586;
        ram[145][63:32] = 32'd2322605034;
        ram[145][95:64] = 32'd3186320755;
        ram[145][127:96] = 32'd2141613643;
        ram[146][31:0] = 32'd4019702194;
        ram[146][63:32] = 32'd1415357636;
        ram[146][95:64] = 32'd3407577517;
        ram[146][127:96] = 32'd976124543;
        ram[147][31:0] = 32'd1568993292;
        ram[147][63:32] = 32'd1522418319;
        ram[147][95:64] = 32'd3186803448;
        ram[147][127:96] = 32'd408415037;
        ram[148][31:0] = 32'd1698532447;
        ram[148][63:32] = 32'd3272624999;
        ram[148][95:64] = 32'd2517975264;
        ram[148][127:96] = 32'd1596839337;
        ram[149][31:0] = 32'd942647997;
        ram[149][63:32] = 32'd2479920114;
        ram[149][95:64] = 32'd4255124355;
        ram[149][127:96] = 32'd982430234;
        ram[150][31:0] = 32'd3556822102;
        ram[150][63:32] = 32'd750890938;
        ram[150][95:64] = 32'd3047685941;
        ram[150][127:96] = 32'd3423135913;
        ram[151][31:0] = 32'd2682490133;
        ram[151][63:32] = 32'd4062492645;
        ram[151][95:64] = 32'd3682415596;
        ram[151][127:96] = 32'd306393857;
        ram[152][31:0] = 32'd1838197034;
        ram[152][63:32] = 32'd412456713;
        ram[152][95:64] = 32'd3240265434;
        ram[152][127:96] = 32'd3431050438;
        ram[153][31:0] = 32'd551188312;
        ram[153][63:32] = 32'd3036714220;
        ram[153][95:64] = 32'd1362451819;
        ram[153][127:96] = 32'd3586907395;
        ram[154][31:0] = 32'd1633853584;
        ram[154][63:32] = 32'd404883268;
        ram[154][95:64] = 32'd172247604;
        ram[154][127:96] = 32'd3850720077;
        ram[155][31:0] = 32'd1355409361;
        ram[155][63:32] = 32'd3559258385;
        ram[155][95:64] = 32'd2576794356;
        ram[155][127:96] = 32'd1096932212;
        ram[156][31:0] = 32'd1317201626;
        ram[156][63:32] = 32'd1251593008;
        ram[156][95:64] = 32'd3713789991;
        ram[156][127:96] = 32'd1679511367;
        ram[157][31:0] = 32'd3449788833;
        ram[157][63:32] = 32'd1317727169;
        ram[157][95:64] = 32'd3548473177;
        ram[157][127:96] = 32'd2390103675;
        ram[158][31:0] = 32'd173501673;
        ram[158][63:32] = 32'd2419434228;
        ram[158][95:64] = 32'd1252027539;
        ram[158][127:96] = 32'd670392651;
        ram[159][31:0] = 32'd130031873;
        ram[159][63:32] = 32'd2435865425;
        ram[159][95:64] = 32'd2854357662;
        ram[159][127:96] = 32'd2378925636;
        ram[160][31:0] = 32'd2328757272;
        ram[160][63:32] = 32'd3611907161;
        ram[160][95:64] = 32'd1175810859;
        ram[160][127:96] = 32'd4248025510;
        ram[161][31:0] = 32'd487448243;
        ram[161][63:32] = 32'd1218724220;
        ram[161][95:64] = 32'd1152709717;
        ram[161][127:96] = 32'd3910443005;
        ram[162][31:0] = 32'd776883759;
        ram[162][63:32] = 32'd3154846827;
        ram[162][95:64] = 32'd1968337716;
        ram[162][127:96] = 32'd2495032494;
        ram[163][31:0] = 32'd1737322648;
        ram[163][63:32] = 32'd726048092;
        ram[163][95:64] = 32'd3127591198;
        ram[163][127:96] = 32'd3509997369;
        ram[164][31:0] = 32'd218457727;
        ram[164][63:32] = 32'd832697036;
        ram[164][95:64] = 32'd420911824;
        ram[164][127:96] = 32'd3715143865;
        ram[165][31:0] = 32'd270341019;
        ram[165][63:32] = 32'd3720845072;
        ram[165][95:64] = 32'd2741441705;
        ram[165][127:96] = 32'd2417445093;
        ram[166][31:0] = 32'd961409848;
        ram[166][63:32] = 32'd1769037600;
        ram[166][95:64] = 32'd3656350260;
        ram[166][127:96] = 32'd2982965549;
        ram[167][31:0] = 32'd3359216141;
        ram[167][63:32] = 32'd420503772;
        ram[167][95:64] = 32'd2483701347;
        ram[167][127:96] = 32'd660543359;
        ram[168][31:0] = 32'd1705980159;
        ram[168][63:32] = 32'd3460743945;
        ram[168][95:64] = 32'd1495437377;
        ram[168][127:96] = 32'd3828766155;
        ram[169][31:0] = 32'd1442188537;
        ram[169][63:32] = 32'd4176733826;
        ram[169][95:64] = 32'd1095345628;
        ram[169][127:96] = 32'd1411385993;
        ram[170][31:0] = 32'd2167949268;
        ram[170][63:32] = 32'd3780431380;
        ram[170][95:64] = 32'd522462869;
        ram[170][127:96] = 32'd452619150;
        ram[171][31:0] = 32'd3800346499;
        ram[171][63:32] = 32'd2566337623;
        ram[171][95:64] = 32'd3310495543;
        ram[171][127:96] = 32'd208276597;
        ram[172][31:0] = 32'd3075220499;
        ram[172][63:32] = 32'd1724620145;
        ram[172][95:64] = 32'd3106437015;
        ram[172][127:96] = 32'd3982442458;
        ram[173][31:0] = 32'd1622816285;
        ram[173][63:32] = 32'd3113725398;
        ram[173][95:64] = 32'd62309893;
        ram[173][127:96] = 32'd2282602147;
        ram[174][31:0] = 32'd274861910;
        ram[174][63:32] = 32'd3794458561;
        ram[174][95:64] = 32'd154010637;
        ram[174][127:96] = 32'd1566213253;
        ram[175][31:0] = 32'd3305228857;
        ram[175][63:32] = 32'd3933897631;
        ram[175][95:64] = 32'd2033116760;
        ram[175][127:96] = 32'd2171400527;
        ram[176][31:0] = 32'd851967156;
        ram[176][63:32] = 32'd1050986732;
        ram[176][95:64] = 32'd1115261743;
        ram[176][127:96] = 32'd2518819451;
        ram[177][31:0] = 32'd3912899891;
        ram[177][63:32] = 32'd224129802;
        ram[177][95:64] = 32'd3528144181;
        ram[177][127:96] = 32'd2022344989;
        ram[178][31:0] = 32'd1962337977;
        ram[178][63:32] = 32'd3785505943;
        ram[178][95:64] = 32'd2379751579;
        ram[178][127:96] = 32'd1410684338;
        ram[179][31:0] = 32'd1756901617;
        ram[179][63:32] = 32'd1559616511;
        ram[179][95:64] = 32'd3058537315;
        ram[179][127:96] = 32'd2098011958;
        ram[180][31:0] = 32'd1279230111;
        ram[180][63:32] = 32'd3305804503;
        ram[180][95:64] = 32'd3177944058;
        ram[180][127:96] = 32'd1900853036;
        ram[181][31:0] = 32'd3326485598;
        ram[181][63:32] = 32'd1069406399;
        ram[181][95:64] = 32'd4007895896;
        ram[181][127:96] = 32'd2861577116;
        ram[182][31:0] = 32'd2130178182;
        ram[182][63:32] = 32'd2078345693;
        ram[182][95:64] = 32'd3961431253;
        ram[182][127:96] = 32'd3189626759;
        ram[183][31:0] = 32'd999882873;
        ram[183][63:32] = 32'd4174718137;
        ram[183][95:64] = 32'd2715359325;
        ram[183][127:96] = 32'd3254548139;
        ram[184][31:0] = 32'd858000912;
        ram[184][63:32] = 32'd2707504632;
        ram[184][95:64] = 32'd2936876441;
        ram[184][127:96] = 32'd452365728;
        ram[185][31:0] = 32'd3202433012;
        ram[185][63:32] = 32'd4113207875;
        ram[185][95:64] = 32'd3275234631;
        ram[185][127:96] = 32'd426086645;
        ram[186][31:0] = 32'd2404663132;
        ram[186][63:32] = 32'd3467710558;
        ram[186][95:64] = 32'd1546724884;
        ram[186][127:96] = 32'd89299359;
        ram[187][31:0] = 32'd740310607;
        ram[187][63:32] = 32'd3249465326;
        ram[187][95:64] = 32'd3873234694;
        ram[187][127:96] = 32'd2207759834;
        ram[188][31:0] = 32'd1797288606;
        ram[188][63:32] = 32'd214909213;
        ram[188][95:64] = 32'd2117224723;
        ram[188][127:96] = 32'd2779572929;
        ram[189][31:0] = 32'd3136622451;
        ram[189][63:32] = 32'd2524440412;
        ram[189][95:64] = 32'd1681383457;
        ram[189][127:96] = 32'd2903484336;
        ram[190][31:0] = 32'd2966775552;
        ram[190][63:32] = 32'd1166682391;
        ram[190][95:64] = 32'd2301973470;
        ram[190][127:96] = 32'd2747999055;
        ram[191][31:0] = 32'd1805789468;
        ram[191][63:32] = 32'd1817152200;
        ram[191][95:64] = 32'd1789751731;
        ram[191][127:96] = 32'd2928940173;
        ram[192][31:0] = 32'd2226595292;
        ram[192][63:32] = 32'd3339946973;
        ram[192][95:64] = 32'd968883625;
        ram[192][127:96] = 32'd1262750963;
        ram[193][31:0] = 32'd4061278725;
        ram[193][63:32] = 32'd4219261467;
        ram[193][95:64] = 32'd877880049;
        ram[193][127:96] = 32'd3939170061;
        ram[194][31:0] = 32'd2515051088;
        ram[194][63:32] = 32'd3175216081;
        ram[194][95:64] = 32'd2576340339;
        ram[194][127:96] = 32'd1916648810;
        ram[195][31:0] = 32'd2476818174;
        ram[195][63:32] = 32'd2253784569;
        ram[195][95:64] = 32'd357526767;
        ram[195][127:96] = 32'd600722239;
        ram[196][31:0] = 32'd560379488;
        ram[196][63:32] = 32'd2691045821;
        ram[196][95:64] = 32'd876002850;
        ram[196][127:96] = 32'd109264237;
        ram[197][31:0] = 32'd1639691474;
        ram[197][63:32] = 32'd2090407313;
        ram[197][95:64] = 32'd1890470687;
        ram[197][127:96] = 32'd496190147;
        ram[198][31:0] = 32'd4118310628;
        ram[198][63:32] = 32'd1132372465;
        ram[198][95:64] = 32'd2371798522;
        ram[198][127:96] = 32'd2253800365;
        ram[199][31:0] = 32'd1668815192;
        ram[199][63:32] = 32'd3852826982;
        ram[199][95:64] = 32'd1995026993;
        ram[199][127:96] = 32'd3803697363;
        ram[200][31:0] = 32'd3694851582;
        ram[200][63:32] = 32'd996574026;
        ram[200][95:64] = 32'd3175044348;
        ram[200][127:96] = 32'd3908749165;
        ram[201][31:0] = 32'd3237418627;
        ram[201][63:32] = 32'd627959300;
        ram[201][95:64] = 32'd3113296974;
        ram[201][127:96] = 32'd1709814211;
        ram[202][31:0] = 32'd3076343433;
        ram[202][63:32] = 32'd1538329166;
        ram[202][95:64] = 32'd914364136;
        ram[202][127:96] = 32'd3314424292;
        ram[203][31:0] = 32'd2940558418;
        ram[203][63:32] = 32'd1334329655;
        ram[203][95:64] = 32'd2882689993;
        ram[203][127:96] = 32'd933026224;
        ram[204][31:0] = 32'd96275483;
        ram[204][63:32] = 32'd1666061305;
        ram[204][95:64] = 32'd160882647;
        ram[204][127:96] = 32'd3916228144;
        ram[205][31:0] = 32'd3676412073;
        ram[205][63:32] = 32'd707615435;
        ram[205][95:64] = 32'd661016934;
        ram[205][127:96] = 32'd4008531324;
        ram[206][31:0] = 32'd397224463;
        ram[206][63:32] = 32'd276834200;
        ram[206][95:64] = 32'd251042263;
        ram[206][127:96] = 32'd494622755;
        ram[207][31:0] = 32'd3353314327;
        ram[207][63:32] = 32'd2221576581;
        ram[207][95:64] = 32'd1059674500;
        ram[207][127:96] = 32'd11545355;
        ram[208][31:0] = 32'd2809961330;
        ram[208][63:32] = 32'd1455017460;
        ram[208][95:64] = 32'd1361242571;
        ram[208][127:96] = 32'd1213873382;
        ram[209][31:0] = 32'd2037704408;
        ram[209][63:32] = 32'd1657911559;
        ram[209][95:64] = 32'd924586107;
        ram[209][127:96] = 32'd1862425237;
        ram[210][31:0] = 32'd3618252464;
        ram[210][63:32] = 32'd209372675;
        ram[210][95:64] = 32'd2607202746;
        ram[210][127:96] = 32'd4105319985;
        ram[211][31:0] = 32'd4108930760;
        ram[211][63:32] = 32'd3010963361;
        ram[211][95:64] = 32'd3871268654;
        ram[211][127:96] = 32'd2811533726;
        ram[212][31:0] = 32'd4074463617;
        ram[212][63:32] = 32'd4029825875;
        ram[212][95:64] = 32'd1441541226;
        ram[212][127:96] = 32'd3497740514;
        ram[213][31:0] = 32'd2241971371;
        ram[213][63:32] = 32'd2928255153;
        ram[213][95:64] = 32'd804645170;
        ram[213][127:96] = 32'd2688237503;
        ram[214][31:0] = 32'd3274644583;
        ram[214][63:32] = 32'd2231454879;
        ram[214][95:64] = 32'd4000613725;
        ram[214][127:96] = 32'd544317971;
        ram[215][31:0] = 32'd3246602886;
        ram[215][63:32] = 32'd1495467381;
        ram[215][95:64] = 32'd3532219985;
        ram[215][127:96] = 32'd2533925369;
        ram[216][31:0] = 32'd385659595;
        ram[216][63:32] = 32'd3491167284;
        ram[216][95:64] = 32'd1790450436;
        ram[216][127:96] = 32'd4125868575;
        ram[217][31:0] = 32'd3743578642;
        ram[217][63:32] = 32'd2026266664;
        ram[217][95:64] = 32'd2235229089;
        ram[217][127:96] = 32'd3307625235;
        ram[218][31:0] = 32'd3804298615;
        ram[218][63:32] = 32'd3342053540;
        ram[218][95:64] = 32'd3793369460;
        ram[218][127:96] = 32'd4043269648;
        ram[219][31:0] = 32'd1362121102;
        ram[219][63:32] = 32'd2198385985;
        ram[219][95:64] = 32'd886953612;
        ram[219][127:96] = 32'd3146529035;
        ram[220][31:0] = 32'd1513837228;
        ram[220][63:32] = 32'd1205481735;
        ram[220][95:64] = 32'd2485169474;
        ram[220][127:96] = 32'd3455419731;
        ram[221][31:0] = 32'd1603698784;
        ram[221][63:32] = 32'd169185942;
        ram[221][95:64] = 32'd3848846976;
        ram[221][127:96] = 32'd2461902253;
        ram[222][31:0] = 32'd2681275051;
        ram[222][63:32] = 32'd2057980656;
        ram[222][95:64] = 32'd1018830267;
        ram[222][127:96] = 32'd4197184161;
        ram[223][31:0] = 32'd1771063249;
        ram[223][63:32] = 32'd2729806528;
        ram[223][95:64] = 32'd1657957379;
        ram[223][127:96] = 32'd1344756801;
        ram[224][31:0] = 32'd1203527177;
        ram[224][63:32] = 32'd1983065030;
        ram[224][95:64] = 32'd4257032184;
        ram[224][127:96] = 32'd2405277136;
        ram[225][31:0] = 32'd3781980178;
        ram[225][63:32] = 32'd467252117;
        ram[225][95:64] = 32'd1936707642;
        ram[225][127:96] = 32'd2261707201;
        ram[226][31:0] = 32'd2619155067;
        ram[226][63:32] = 32'd866381383;
        ram[226][95:64] = 32'd1994273950;
        ram[226][127:96] = 32'd1385986733;
        ram[227][31:0] = 32'd214893740;
        ram[227][63:32] = 32'd3200669720;
        ram[227][95:64] = 32'd2791318259;
        ram[227][127:96] = 32'd360531280;
        ram[228][31:0] = 32'd1323603140;
        ram[228][63:32] = 32'd1701002144;
        ram[228][95:64] = 32'd617611722;
        ram[228][127:96] = 32'd316048180;
        ram[229][31:0] = 32'd2296523743;
        ram[229][63:32] = 32'd347883434;
        ram[229][95:64] = 32'd1901704297;
        ram[229][127:96] = 32'd1993211956;
        ram[230][31:0] = 32'd1049468648;
        ram[230][63:32] = 32'd1768926262;
        ram[230][95:64] = 32'd268862713;
        ram[230][127:96] = 32'd2554414221;
        ram[231][31:0] = 32'd2196417372;
        ram[231][63:32] = 32'd74622926;
        ram[231][95:64] = 32'd2262293352;
        ram[231][127:96] = 32'd3488619352;
        ram[232][31:0] = 32'd3420167902;
        ram[232][63:32] = 32'd940344392;
        ram[232][95:64] = 32'd1966535596;
        ram[232][127:96] = 32'd3103550827;
        ram[233][31:0] = 32'd2930470201;
        ram[233][63:32] = 32'd2511644972;
        ram[233][95:64] = 32'd2823866363;
        ram[233][127:96] = 32'd1717104902;
        ram[234][31:0] = 32'd3123676491;
        ram[234][63:32] = 32'd2203028531;
        ram[234][95:64] = 32'd2400356313;
        ram[234][127:96] = 32'd2075534042;
        ram[235][31:0] = 32'd1707455229;
        ram[235][63:32] = 32'd2844599084;
        ram[235][95:64] = 32'd857066257;
        ram[235][127:96] = 32'd3573192684;
        ram[236][31:0] = 32'd1106836672;
        ram[236][63:32] = 32'd4038263291;
        ram[236][95:64] = 32'd3719653609;
        ram[236][127:96] = 32'd3478032258;
        ram[237][31:0] = 32'd1347233679;
        ram[237][63:32] = 32'd318477808;
        ram[237][95:64] = 32'd1837511223;
        ram[237][127:96] = 32'd1276682534;
        ram[238][31:0] = 32'd3841582932;
        ram[238][63:32] = 32'd1358315614;
        ram[238][95:64] = 32'd3948916793;
        ram[238][127:96] = 32'd976392251;
        ram[239][31:0] = 32'd604891091;
        ram[239][63:32] = 32'd2766494036;
        ram[239][95:64] = 32'd3933242076;
        ram[239][127:96] = 32'd1529856229;
        ram[240][31:0] = 32'd1948195766;
        ram[240][63:32] = 32'd2424908381;
        ram[240][95:64] = 32'd1061798646;
        ram[240][127:96] = 32'd116665739;
        ram[241][31:0] = 32'd864540540;
        ram[241][63:32] = 32'd3248282811;
        ram[241][95:64] = 32'd4155125915;
        ram[241][127:96] = 32'd2231060372;
        ram[242][31:0] = 32'd1749865633;
        ram[242][63:32] = 32'd2080802869;
        ram[242][95:64] = 32'd2451347637;
        ram[242][127:96] = 32'd713104100;
        ram[243][31:0] = 32'd3792588729;
        ram[243][63:32] = 32'd1940515451;
        ram[243][95:64] = 32'd947401983;
        ram[243][127:96] = 32'd3022759963;
        ram[244][31:0] = 32'd3450979905;
        ram[244][63:32] = 32'd3853008963;
        ram[244][95:64] = 32'd505129006;
        ram[244][127:96] = 32'd3351282188;
        ram[245][31:0] = 32'd127768736;
        ram[245][63:32] = 32'd1414503463;
        ram[245][95:64] = 32'd681903484;
        ram[245][127:96] = 32'd1650122225;
        ram[246][31:0] = 32'd2979938981;
        ram[246][63:32] = 32'd2125246417;
        ram[246][95:64] = 32'd2058768324;
        ram[246][127:96] = 32'd2669326286;
        ram[247][31:0] = 32'd1629806814;
        ram[247][63:32] = 32'd867504778;
        ram[247][95:64] = 32'd4133797271;
        ram[247][127:96] = 32'd4151446151;
        ram[248][31:0] = 32'd112184677;
        ram[248][63:32] = 32'd3829262925;
        ram[248][95:64] = 32'd3294305116;
        ram[248][127:96] = 32'd1145317896;
        ram[249][31:0] = 32'd428556190;
        ram[249][63:32] = 32'd3032800360;
        ram[249][95:64] = 32'd4049855863;
        ram[249][127:96] = 32'd3909732291;
        ram[250][31:0] = 32'd3487038663;
        ram[250][63:32] = 32'd3081669374;
        ram[250][95:64] = 32'd587228443;
        ram[250][127:96] = 32'd3486094991;
        ram[251][31:0] = 32'd3494997726;
        ram[251][63:32] = 32'd2647342235;
        ram[251][95:64] = 32'd4197983772;
        ram[251][127:96] = 32'd492031920;
        ram[252][31:0] = 32'd2946475741;
        ram[252][63:32] = 32'd994495003;
        ram[252][95:64] = 32'd704857744;
        ram[252][127:96] = 32'd359423007;
        ram[253][31:0] = 32'd3811102047;
        ram[253][63:32] = 32'd2547033048;
        ram[253][95:64] = 32'd1358387716;
        ram[253][127:96] = 32'd2574971247;
        ram[254][31:0] = 32'd3018854002;
        ram[254][63:32] = 32'd4080120458;
        ram[254][95:64] = 32'd4106663678;
        ram[254][127:96] = 32'd2406923194;
        ram[255][31:0] = 32'd2038773800;
        ram[255][63:32] = 32'd1031762782;
        ram[255][95:64] = 32'd1277705246;
        ram[255][127:96] = 32'd2086004592;

    end
    always @(posedge clk) begin
        addr_r <= raddr;
        if(we) ram[waddr] <= din;
    end
    assign dout = ram[addr_r]; 

endmodule
